// Generator : SpinalHDL v1.9.4    git head : 270018552577f3bb8e5339ee2583c9c22d324215
// Component : uSystolicArray
// Git hash  : 95d4b99c2c5c0c9e41b84111df30141758565e63

`timescale 1ns/1ps

module uSystolicArray (
  input  wire [15:0]   io_enable_i,
  input  wire [15:0]   io_clear_i,
  input  wire [15:0]   io_mac_done,
  input  wire [15:0]   io_enable_w,
  input  wire [15:0]   io_clear_w,
  input  wire [15:0]   io_enable_o,
  input  wire [15:0]   io_clear_o,
  input  wire [15:0]   io_ifm_0,
  input  wire [15:0]   io_ifm_1,
  input  wire [15:0]   io_ifm_2,
  input  wire [15:0]   io_ifm_3,
  input  wire [15:0]   io_ifm_4,
  input  wire [15:0]   io_ifm_5,
  input  wire [15:0]   io_ifm_6,
  input  wire [15:0]   io_ifm_7,
  input  wire [15:0]   io_ifm_8,
  input  wire [15:0]   io_ifm_9,
  input  wire [15:0]   io_ifm_10,
  input  wire [15:0]   io_ifm_11,
  input  wire [15:0]   io_ifm_12,
  input  wire [15:0]   io_ifm_13,
  input  wire [15:0]   io_ifm_14,
  input  wire [15:0]   io_ifm_15,
  input  wire [15:0]   io_wght_sign,
  input  wire [14:0]   io_wght_abs_0,
  input  wire [14:0]   io_wght_abs_1,
  input  wire [14:0]   io_wght_abs_2,
  input  wire [14:0]   io_wght_abs_3,
  input  wire [14:0]   io_wght_abs_4,
  input  wire [14:0]   io_wght_abs_5,
  input  wire [14:0]   io_wght_abs_6,
  input  wire [14:0]   io_wght_abs_7,
  input  wire [14:0]   io_wght_abs_8,
  input  wire [14:0]   io_wght_abs_9,
  input  wire [14:0]   io_wght_abs_10,
  input  wire [14:0]   io_wght_abs_11,
  input  wire [14:0]   io_wght_abs_12,
  input  wire [14:0]   io_wght_abs_13,
  input  wire [14:0]   io_wght_abs_14,
  input  wire [14:0]   io_wght_abs_15,
  output wire [31:0]   io_ofm_0,
  output wire [31:0]   io_ofm_1,
  output wire [31:0]   io_ofm_2,
  output wire [31:0]   io_ofm_3,
  output wire [31:0]   io_ofm_4,
  output wire [31:0]   io_ofm_5,
  output wire [31:0]   io_ofm_6,
  output wire [31:0]   io_ofm_7,
  output wire [31:0]   io_ofm_8,
  output wire [31:0]   io_ofm_9,
  output wire [31:0]   io_ofm_10,
  output wire [31:0]   io_ofm_11,
  output wire [31:0]   io_ofm_12,
  output wire [31:0]   io_ofm_13,
  output wire [31:0]   io_ofm_14,
  output wire [31:0]   io_ofm_15,
  input  wire          clk,
  input  wire          reset
);

  wire                uSystolicPEBorder_16_io_mac_done;
  wire                uSystolicPEBorder_16_io_enable_i;
  wire                uSystolicPEBorder_16_io_clear_i;
  wire                uSystolicPEBorder_16_io_enable_w;
  wire                uSystolicPEBorder_16_io_clear_w;
  wire                uSystolicPEBorder_16_io_enable_o;
  wire                uSystolicPEBorder_16_io_clear_o;
  wire                uSystolicPE_240_io_mac_done;
  wire                uSystolicPE_240_io_enable_i;
  wire                uSystolicPE_240_io_clear_i;
  wire                uSystolicPE_240_io_enable_w;
  wire                uSystolicPE_240_io_clear_w;
  wire                uSystolicPE_240_io_enable_o;
  wire                uSystolicPE_240_io_clear_o;
  wire                uSystolicPE_241_io_mac_done;
  wire                uSystolicPE_241_io_enable_i;
  wire                uSystolicPE_241_io_clear_i;
  wire                uSystolicPE_241_io_enable_w;
  wire                uSystolicPE_241_io_clear_w;
  wire                uSystolicPE_241_io_enable_o;
  wire                uSystolicPE_241_io_clear_o;
  wire                uSystolicPE_242_io_mac_done;
  wire                uSystolicPE_242_io_enable_i;
  wire                uSystolicPE_242_io_clear_i;
  wire                uSystolicPE_242_io_enable_w;
  wire                uSystolicPE_242_io_clear_w;
  wire                uSystolicPE_242_io_enable_o;
  wire                uSystolicPE_242_io_clear_o;
  wire                uSystolicPE_243_io_mac_done;
  wire                uSystolicPE_243_io_enable_i;
  wire                uSystolicPE_243_io_clear_i;
  wire                uSystolicPE_243_io_enable_w;
  wire                uSystolicPE_243_io_clear_w;
  wire                uSystolicPE_243_io_enable_o;
  wire                uSystolicPE_243_io_clear_o;
  wire                uSystolicPE_244_io_mac_done;
  wire                uSystolicPE_244_io_enable_i;
  wire                uSystolicPE_244_io_clear_i;
  wire                uSystolicPE_244_io_enable_w;
  wire                uSystolicPE_244_io_clear_w;
  wire                uSystolicPE_244_io_enable_o;
  wire                uSystolicPE_244_io_clear_o;
  wire                uSystolicPE_245_io_mac_done;
  wire                uSystolicPE_245_io_enable_i;
  wire                uSystolicPE_245_io_clear_i;
  wire                uSystolicPE_245_io_enable_w;
  wire                uSystolicPE_245_io_clear_w;
  wire                uSystolicPE_245_io_enable_o;
  wire                uSystolicPE_245_io_clear_o;
  wire                uSystolicPE_246_io_mac_done;
  wire                uSystolicPE_246_io_enable_i;
  wire                uSystolicPE_246_io_clear_i;
  wire                uSystolicPE_246_io_enable_w;
  wire                uSystolicPE_246_io_clear_w;
  wire                uSystolicPE_246_io_enable_o;
  wire                uSystolicPE_246_io_clear_o;
  wire                uSystolicPE_247_io_mac_done;
  wire                uSystolicPE_247_io_enable_i;
  wire                uSystolicPE_247_io_clear_i;
  wire                uSystolicPE_247_io_enable_w;
  wire                uSystolicPE_247_io_clear_w;
  wire                uSystolicPE_247_io_enable_o;
  wire                uSystolicPE_247_io_clear_o;
  wire                uSystolicPE_248_io_mac_done;
  wire                uSystolicPE_248_io_enable_i;
  wire                uSystolicPE_248_io_clear_i;
  wire                uSystolicPE_248_io_enable_w;
  wire                uSystolicPE_248_io_clear_w;
  wire                uSystolicPE_248_io_enable_o;
  wire                uSystolicPE_248_io_clear_o;
  wire                uSystolicPE_249_io_mac_done;
  wire                uSystolicPE_249_io_enable_i;
  wire                uSystolicPE_249_io_clear_i;
  wire                uSystolicPE_249_io_enable_w;
  wire                uSystolicPE_249_io_clear_w;
  wire                uSystolicPE_249_io_enable_o;
  wire                uSystolicPE_249_io_clear_o;
  wire                uSystolicPE_250_io_mac_done;
  wire                uSystolicPE_250_io_enable_i;
  wire                uSystolicPE_250_io_clear_i;
  wire                uSystolicPE_250_io_enable_w;
  wire                uSystolicPE_250_io_clear_w;
  wire                uSystolicPE_250_io_enable_o;
  wire                uSystolicPE_250_io_clear_o;
  wire                uSystolicPE_251_io_mac_done;
  wire                uSystolicPE_251_io_enable_i;
  wire                uSystolicPE_251_io_clear_i;
  wire                uSystolicPE_251_io_enable_w;
  wire                uSystolicPE_251_io_clear_w;
  wire                uSystolicPE_251_io_enable_o;
  wire                uSystolicPE_251_io_clear_o;
  wire                uSystolicPE_252_io_mac_done;
  wire                uSystolicPE_252_io_enable_i;
  wire                uSystolicPE_252_io_clear_i;
  wire                uSystolicPE_252_io_enable_w;
  wire                uSystolicPE_252_io_clear_w;
  wire                uSystolicPE_252_io_enable_o;
  wire                uSystolicPE_252_io_clear_o;
  wire                uSystolicPE_253_io_mac_done;
  wire                uSystolicPE_253_io_enable_i;
  wire                uSystolicPE_253_io_clear_i;
  wire                uSystolicPE_253_io_enable_w;
  wire                uSystolicPE_253_io_clear_w;
  wire                uSystolicPE_253_io_enable_o;
  wire                uSystolicPE_253_io_clear_o;
  wire                uSystolicPE_254_io_mac_done;
  wire                uSystolicPE_254_io_enable_i;
  wire                uSystolicPE_254_io_clear_i;
  wire                uSystolicPE_254_io_enable_w;
  wire                uSystolicPE_254_io_clear_w;
  wire                uSystolicPE_254_io_enable_o;
  wire                uSystolicPE_254_io_clear_o;
  wire                uSystolicPEBorder_17_io_mac_done;
  wire                uSystolicPEBorder_17_io_enable_i;
  wire                uSystolicPEBorder_17_io_clear_i;
  wire                uSystolicPEBorder_17_io_enable_w;
  wire                uSystolicPEBorder_17_io_clear_w;
  wire                uSystolicPEBorder_17_io_enable_o;
  wire                uSystolicPEBorder_17_io_clear_o;
  wire                uSystolicPE_255_io_mac_done;
  wire                uSystolicPE_255_io_enable_i;
  wire                uSystolicPE_255_io_clear_i;
  wire                uSystolicPE_255_io_enable_w;
  wire                uSystolicPE_255_io_clear_w;
  wire                uSystolicPE_255_io_enable_o;
  wire                uSystolicPE_255_io_clear_o;
  wire                uSystolicPE_256_io_mac_done;
  wire                uSystolicPE_256_io_enable_i;
  wire                uSystolicPE_256_io_clear_i;
  wire                uSystolicPE_256_io_enable_w;
  wire                uSystolicPE_256_io_clear_w;
  wire                uSystolicPE_256_io_enable_o;
  wire                uSystolicPE_256_io_clear_o;
  wire                uSystolicPE_257_io_mac_done;
  wire                uSystolicPE_257_io_enable_i;
  wire                uSystolicPE_257_io_clear_i;
  wire                uSystolicPE_257_io_enable_w;
  wire                uSystolicPE_257_io_clear_w;
  wire                uSystolicPE_257_io_enable_o;
  wire                uSystolicPE_257_io_clear_o;
  wire                uSystolicPE_258_io_mac_done;
  wire                uSystolicPE_258_io_enable_i;
  wire                uSystolicPE_258_io_clear_i;
  wire                uSystolicPE_258_io_enable_w;
  wire                uSystolicPE_258_io_clear_w;
  wire                uSystolicPE_258_io_enable_o;
  wire                uSystolicPE_258_io_clear_o;
  wire                uSystolicPE_259_io_mac_done;
  wire                uSystolicPE_259_io_enable_i;
  wire                uSystolicPE_259_io_clear_i;
  wire                uSystolicPE_259_io_enable_w;
  wire                uSystolicPE_259_io_clear_w;
  wire                uSystolicPE_259_io_enable_o;
  wire                uSystolicPE_259_io_clear_o;
  wire                uSystolicPE_260_io_mac_done;
  wire                uSystolicPE_260_io_enable_i;
  wire                uSystolicPE_260_io_clear_i;
  wire                uSystolicPE_260_io_enable_w;
  wire                uSystolicPE_260_io_clear_w;
  wire                uSystolicPE_260_io_enable_o;
  wire                uSystolicPE_260_io_clear_o;
  wire                uSystolicPE_261_io_mac_done;
  wire                uSystolicPE_261_io_enable_i;
  wire                uSystolicPE_261_io_clear_i;
  wire                uSystolicPE_261_io_enable_w;
  wire                uSystolicPE_261_io_clear_w;
  wire                uSystolicPE_261_io_enable_o;
  wire                uSystolicPE_261_io_clear_o;
  wire                uSystolicPE_262_io_mac_done;
  wire                uSystolicPE_262_io_enable_i;
  wire                uSystolicPE_262_io_clear_i;
  wire                uSystolicPE_262_io_enable_w;
  wire                uSystolicPE_262_io_clear_w;
  wire                uSystolicPE_262_io_enable_o;
  wire                uSystolicPE_262_io_clear_o;
  wire                uSystolicPE_263_io_mac_done;
  wire                uSystolicPE_263_io_enable_i;
  wire                uSystolicPE_263_io_clear_i;
  wire                uSystolicPE_263_io_enable_w;
  wire                uSystolicPE_263_io_clear_w;
  wire                uSystolicPE_263_io_enable_o;
  wire                uSystolicPE_263_io_clear_o;
  wire                uSystolicPE_264_io_mac_done;
  wire                uSystolicPE_264_io_enable_i;
  wire                uSystolicPE_264_io_clear_i;
  wire                uSystolicPE_264_io_enable_w;
  wire                uSystolicPE_264_io_clear_w;
  wire                uSystolicPE_264_io_enable_o;
  wire                uSystolicPE_264_io_clear_o;
  wire                uSystolicPE_265_io_mac_done;
  wire                uSystolicPE_265_io_enable_i;
  wire                uSystolicPE_265_io_clear_i;
  wire                uSystolicPE_265_io_enable_w;
  wire                uSystolicPE_265_io_clear_w;
  wire                uSystolicPE_265_io_enable_o;
  wire                uSystolicPE_265_io_clear_o;
  wire                uSystolicPE_266_io_mac_done;
  wire                uSystolicPE_266_io_enable_i;
  wire                uSystolicPE_266_io_clear_i;
  wire                uSystolicPE_266_io_enable_w;
  wire                uSystolicPE_266_io_clear_w;
  wire                uSystolicPE_266_io_enable_o;
  wire                uSystolicPE_266_io_clear_o;
  wire                uSystolicPE_267_io_mac_done;
  wire                uSystolicPE_267_io_enable_i;
  wire                uSystolicPE_267_io_clear_i;
  wire                uSystolicPE_267_io_enable_w;
  wire                uSystolicPE_267_io_clear_w;
  wire                uSystolicPE_267_io_enable_o;
  wire                uSystolicPE_267_io_clear_o;
  wire                uSystolicPE_268_io_mac_done;
  wire                uSystolicPE_268_io_enable_i;
  wire                uSystolicPE_268_io_clear_i;
  wire                uSystolicPE_268_io_enable_w;
  wire                uSystolicPE_268_io_clear_w;
  wire                uSystolicPE_268_io_enable_o;
  wire                uSystolicPE_268_io_clear_o;
  wire                uSystolicPE_269_io_mac_done;
  wire                uSystolicPE_269_io_enable_i;
  wire                uSystolicPE_269_io_clear_i;
  wire                uSystolicPE_269_io_enable_w;
  wire                uSystolicPE_269_io_clear_w;
  wire                uSystolicPE_269_io_enable_o;
  wire                uSystolicPE_269_io_clear_o;
  wire                uSystolicPEBorder_18_io_mac_done;
  wire                uSystolicPEBorder_18_io_enable_i;
  wire                uSystolicPEBorder_18_io_clear_i;
  wire                uSystolicPEBorder_18_io_enable_w;
  wire                uSystolicPEBorder_18_io_clear_w;
  wire                uSystolicPEBorder_18_io_enable_o;
  wire                uSystolicPEBorder_18_io_clear_o;
  wire                uSystolicPE_270_io_mac_done;
  wire                uSystolicPE_270_io_enable_i;
  wire                uSystolicPE_270_io_clear_i;
  wire                uSystolicPE_270_io_enable_w;
  wire                uSystolicPE_270_io_clear_w;
  wire                uSystolicPE_270_io_enable_o;
  wire                uSystolicPE_270_io_clear_o;
  wire                uSystolicPE_271_io_mac_done;
  wire                uSystolicPE_271_io_enable_i;
  wire                uSystolicPE_271_io_clear_i;
  wire                uSystolicPE_271_io_enable_w;
  wire                uSystolicPE_271_io_clear_w;
  wire                uSystolicPE_271_io_enable_o;
  wire                uSystolicPE_271_io_clear_o;
  wire                uSystolicPE_272_io_mac_done;
  wire                uSystolicPE_272_io_enable_i;
  wire                uSystolicPE_272_io_clear_i;
  wire                uSystolicPE_272_io_enable_w;
  wire                uSystolicPE_272_io_clear_w;
  wire                uSystolicPE_272_io_enable_o;
  wire                uSystolicPE_272_io_clear_o;
  wire                uSystolicPE_273_io_mac_done;
  wire                uSystolicPE_273_io_enable_i;
  wire                uSystolicPE_273_io_clear_i;
  wire                uSystolicPE_273_io_enable_w;
  wire                uSystolicPE_273_io_clear_w;
  wire                uSystolicPE_273_io_enable_o;
  wire                uSystolicPE_273_io_clear_o;
  wire                uSystolicPE_274_io_mac_done;
  wire                uSystolicPE_274_io_enable_i;
  wire                uSystolicPE_274_io_clear_i;
  wire                uSystolicPE_274_io_enable_w;
  wire                uSystolicPE_274_io_clear_w;
  wire                uSystolicPE_274_io_enable_o;
  wire                uSystolicPE_274_io_clear_o;
  wire                uSystolicPE_275_io_mac_done;
  wire                uSystolicPE_275_io_enable_i;
  wire                uSystolicPE_275_io_clear_i;
  wire                uSystolicPE_275_io_enable_w;
  wire                uSystolicPE_275_io_clear_w;
  wire                uSystolicPE_275_io_enable_o;
  wire                uSystolicPE_275_io_clear_o;
  wire                uSystolicPE_276_io_mac_done;
  wire                uSystolicPE_276_io_enable_i;
  wire                uSystolicPE_276_io_clear_i;
  wire                uSystolicPE_276_io_enable_w;
  wire                uSystolicPE_276_io_clear_w;
  wire                uSystolicPE_276_io_enable_o;
  wire                uSystolicPE_276_io_clear_o;
  wire                uSystolicPE_277_io_mac_done;
  wire                uSystolicPE_277_io_enable_i;
  wire                uSystolicPE_277_io_clear_i;
  wire                uSystolicPE_277_io_enable_w;
  wire                uSystolicPE_277_io_clear_w;
  wire                uSystolicPE_277_io_enable_o;
  wire                uSystolicPE_277_io_clear_o;
  wire                uSystolicPE_278_io_mac_done;
  wire                uSystolicPE_278_io_enable_i;
  wire                uSystolicPE_278_io_clear_i;
  wire                uSystolicPE_278_io_enable_w;
  wire                uSystolicPE_278_io_clear_w;
  wire                uSystolicPE_278_io_enable_o;
  wire                uSystolicPE_278_io_clear_o;
  wire                uSystolicPE_279_io_mac_done;
  wire                uSystolicPE_279_io_enable_i;
  wire                uSystolicPE_279_io_clear_i;
  wire                uSystolicPE_279_io_enable_w;
  wire                uSystolicPE_279_io_clear_w;
  wire                uSystolicPE_279_io_enable_o;
  wire                uSystolicPE_279_io_clear_o;
  wire                uSystolicPE_280_io_mac_done;
  wire                uSystolicPE_280_io_enable_i;
  wire                uSystolicPE_280_io_clear_i;
  wire                uSystolicPE_280_io_enable_w;
  wire                uSystolicPE_280_io_clear_w;
  wire                uSystolicPE_280_io_enable_o;
  wire                uSystolicPE_280_io_clear_o;
  wire                uSystolicPE_281_io_mac_done;
  wire                uSystolicPE_281_io_enable_i;
  wire                uSystolicPE_281_io_clear_i;
  wire                uSystolicPE_281_io_enable_w;
  wire                uSystolicPE_281_io_clear_w;
  wire                uSystolicPE_281_io_enable_o;
  wire                uSystolicPE_281_io_clear_o;
  wire                uSystolicPE_282_io_mac_done;
  wire                uSystolicPE_282_io_enable_i;
  wire                uSystolicPE_282_io_clear_i;
  wire                uSystolicPE_282_io_enable_w;
  wire                uSystolicPE_282_io_clear_w;
  wire                uSystolicPE_282_io_enable_o;
  wire                uSystolicPE_282_io_clear_o;
  wire                uSystolicPE_283_io_mac_done;
  wire                uSystolicPE_283_io_enable_i;
  wire                uSystolicPE_283_io_clear_i;
  wire                uSystolicPE_283_io_enable_w;
  wire                uSystolicPE_283_io_clear_w;
  wire                uSystolicPE_283_io_enable_o;
  wire                uSystolicPE_283_io_clear_o;
  wire                uSystolicPE_284_io_mac_done;
  wire                uSystolicPE_284_io_enable_i;
  wire                uSystolicPE_284_io_clear_i;
  wire                uSystolicPE_284_io_enable_w;
  wire                uSystolicPE_284_io_clear_w;
  wire                uSystolicPE_284_io_enable_o;
  wire                uSystolicPE_284_io_clear_o;
  wire                uSystolicPEBorder_19_io_mac_done;
  wire                uSystolicPEBorder_19_io_enable_i;
  wire                uSystolicPEBorder_19_io_clear_i;
  wire                uSystolicPEBorder_19_io_enable_w;
  wire                uSystolicPEBorder_19_io_clear_w;
  wire                uSystolicPEBorder_19_io_enable_o;
  wire                uSystolicPEBorder_19_io_clear_o;
  wire                uSystolicPE_285_io_mac_done;
  wire                uSystolicPE_285_io_enable_i;
  wire                uSystolicPE_285_io_clear_i;
  wire                uSystolicPE_285_io_enable_w;
  wire                uSystolicPE_285_io_clear_w;
  wire                uSystolicPE_285_io_enable_o;
  wire                uSystolicPE_285_io_clear_o;
  wire                uSystolicPE_286_io_mac_done;
  wire                uSystolicPE_286_io_enable_i;
  wire                uSystolicPE_286_io_clear_i;
  wire                uSystolicPE_286_io_enable_w;
  wire                uSystolicPE_286_io_clear_w;
  wire                uSystolicPE_286_io_enable_o;
  wire                uSystolicPE_286_io_clear_o;
  wire                uSystolicPE_287_io_mac_done;
  wire                uSystolicPE_287_io_enable_i;
  wire                uSystolicPE_287_io_clear_i;
  wire                uSystolicPE_287_io_enable_w;
  wire                uSystolicPE_287_io_clear_w;
  wire                uSystolicPE_287_io_enable_o;
  wire                uSystolicPE_287_io_clear_o;
  wire                uSystolicPE_288_io_mac_done;
  wire                uSystolicPE_288_io_enable_i;
  wire                uSystolicPE_288_io_clear_i;
  wire                uSystolicPE_288_io_enable_w;
  wire                uSystolicPE_288_io_clear_w;
  wire                uSystolicPE_288_io_enable_o;
  wire                uSystolicPE_288_io_clear_o;
  wire                uSystolicPE_289_io_mac_done;
  wire                uSystolicPE_289_io_enable_i;
  wire                uSystolicPE_289_io_clear_i;
  wire                uSystolicPE_289_io_enable_w;
  wire                uSystolicPE_289_io_clear_w;
  wire                uSystolicPE_289_io_enable_o;
  wire                uSystolicPE_289_io_clear_o;
  wire                uSystolicPE_290_io_mac_done;
  wire                uSystolicPE_290_io_enable_i;
  wire                uSystolicPE_290_io_clear_i;
  wire                uSystolicPE_290_io_enable_w;
  wire                uSystolicPE_290_io_clear_w;
  wire                uSystolicPE_290_io_enable_o;
  wire                uSystolicPE_290_io_clear_o;
  wire                uSystolicPE_291_io_mac_done;
  wire                uSystolicPE_291_io_enable_i;
  wire                uSystolicPE_291_io_clear_i;
  wire                uSystolicPE_291_io_enable_w;
  wire                uSystolicPE_291_io_clear_w;
  wire                uSystolicPE_291_io_enable_o;
  wire                uSystolicPE_291_io_clear_o;
  wire                uSystolicPE_292_io_mac_done;
  wire                uSystolicPE_292_io_enable_i;
  wire                uSystolicPE_292_io_clear_i;
  wire                uSystolicPE_292_io_enable_w;
  wire                uSystolicPE_292_io_clear_w;
  wire                uSystolicPE_292_io_enable_o;
  wire                uSystolicPE_292_io_clear_o;
  wire                uSystolicPE_293_io_mac_done;
  wire                uSystolicPE_293_io_enable_i;
  wire                uSystolicPE_293_io_clear_i;
  wire                uSystolicPE_293_io_enable_w;
  wire                uSystolicPE_293_io_clear_w;
  wire                uSystolicPE_293_io_enable_o;
  wire                uSystolicPE_293_io_clear_o;
  wire                uSystolicPE_294_io_mac_done;
  wire                uSystolicPE_294_io_enable_i;
  wire                uSystolicPE_294_io_clear_i;
  wire                uSystolicPE_294_io_enable_w;
  wire                uSystolicPE_294_io_clear_w;
  wire                uSystolicPE_294_io_enable_o;
  wire                uSystolicPE_294_io_clear_o;
  wire                uSystolicPE_295_io_mac_done;
  wire                uSystolicPE_295_io_enable_i;
  wire                uSystolicPE_295_io_clear_i;
  wire                uSystolicPE_295_io_enable_w;
  wire                uSystolicPE_295_io_clear_w;
  wire                uSystolicPE_295_io_enable_o;
  wire                uSystolicPE_295_io_clear_o;
  wire                uSystolicPE_296_io_mac_done;
  wire                uSystolicPE_296_io_enable_i;
  wire                uSystolicPE_296_io_clear_i;
  wire                uSystolicPE_296_io_enable_w;
  wire                uSystolicPE_296_io_clear_w;
  wire                uSystolicPE_296_io_enable_o;
  wire                uSystolicPE_296_io_clear_o;
  wire                uSystolicPE_297_io_mac_done;
  wire                uSystolicPE_297_io_enable_i;
  wire                uSystolicPE_297_io_clear_i;
  wire                uSystolicPE_297_io_enable_w;
  wire                uSystolicPE_297_io_clear_w;
  wire                uSystolicPE_297_io_enable_o;
  wire                uSystolicPE_297_io_clear_o;
  wire                uSystolicPE_298_io_mac_done;
  wire                uSystolicPE_298_io_enable_i;
  wire                uSystolicPE_298_io_clear_i;
  wire                uSystolicPE_298_io_enable_w;
  wire                uSystolicPE_298_io_clear_w;
  wire                uSystolicPE_298_io_enable_o;
  wire                uSystolicPE_298_io_clear_o;
  wire                uSystolicPE_299_io_mac_done;
  wire                uSystolicPE_299_io_enable_i;
  wire                uSystolicPE_299_io_clear_i;
  wire                uSystolicPE_299_io_enable_w;
  wire                uSystolicPE_299_io_clear_w;
  wire                uSystolicPE_299_io_enable_o;
  wire                uSystolicPE_299_io_clear_o;
  wire                uSystolicPEBorder_20_io_mac_done;
  wire                uSystolicPEBorder_20_io_enable_i;
  wire                uSystolicPEBorder_20_io_clear_i;
  wire                uSystolicPEBorder_20_io_enable_w;
  wire                uSystolicPEBorder_20_io_clear_w;
  wire                uSystolicPEBorder_20_io_enable_o;
  wire                uSystolicPEBorder_20_io_clear_o;
  wire                uSystolicPE_300_io_mac_done;
  wire                uSystolicPE_300_io_enable_i;
  wire                uSystolicPE_300_io_clear_i;
  wire                uSystolicPE_300_io_enable_w;
  wire                uSystolicPE_300_io_clear_w;
  wire                uSystolicPE_300_io_enable_o;
  wire                uSystolicPE_300_io_clear_o;
  wire                uSystolicPE_301_io_mac_done;
  wire                uSystolicPE_301_io_enable_i;
  wire                uSystolicPE_301_io_clear_i;
  wire                uSystolicPE_301_io_enable_w;
  wire                uSystolicPE_301_io_clear_w;
  wire                uSystolicPE_301_io_enable_o;
  wire                uSystolicPE_301_io_clear_o;
  wire                uSystolicPE_302_io_mac_done;
  wire                uSystolicPE_302_io_enable_i;
  wire                uSystolicPE_302_io_clear_i;
  wire                uSystolicPE_302_io_enable_w;
  wire                uSystolicPE_302_io_clear_w;
  wire                uSystolicPE_302_io_enable_o;
  wire                uSystolicPE_302_io_clear_o;
  wire                uSystolicPE_303_io_mac_done;
  wire                uSystolicPE_303_io_enable_i;
  wire                uSystolicPE_303_io_clear_i;
  wire                uSystolicPE_303_io_enable_w;
  wire                uSystolicPE_303_io_clear_w;
  wire                uSystolicPE_303_io_enable_o;
  wire                uSystolicPE_303_io_clear_o;
  wire                uSystolicPE_304_io_mac_done;
  wire                uSystolicPE_304_io_enable_i;
  wire                uSystolicPE_304_io_clear_i;
  wire                uSystolicPE_304_io_enable_w;
  wire                uSystolicPE_304_io_clear_w;
  wire                uSystolicPE_304_io_enable_o;
  wire                uSystolicPE_304_io_clear_o;
  wire                uSystolicPE_305_io_mac_done;
  wire                uSystolicPE_305_io_enable_i;
  wire                uSystolicPE_305_io_clear_i;
  wire                uSystolicPE_305_io_enable_w;
  wire                uSystolicPE_305_io_clear_w;
  wire                uSystolicPE_305_io_enable_o;
  wire                uSystolicPE_305_io_clear_o;
  wire                uSystolicPE_306_io_mac_done;
  wire                uSystolicPE_306_io_enable_i;
  wire                uSystolicPE_306_io_clear_i;
  wire                uSystolicPE_306_io_enable_w;
  wire                uSystolicPE_306_io_clear_w;
  wire                uSystolicPE_306_io_enable_o;
  wire                uSystolicPE_306_io_clear_o;
  wire                uSystolicPE_307_io_mac_done;
  wire                uSystolicPE_307_io_enable_i;
  wire                uSystolicPE_307_io_clear_i;
  wire                uSystolicPE_307_io_enable_w;
  wire                uSystolicPE_307_io_clear_w;
  wire                uSystolicPE_307_io_enable_o;
  wire                uSystolicPE_307_io_clear_o;
  wire                uSystolicPE_308_io_mac_done;
  wire                uSystolicPE_308_io_enable_i;
  wire                uSystolicPE_308_io_clear_i;
  wire                uSystolicPE_308_io_enable_w;
  wire                uSystolicPE_308_io_clear_w;
  wire                uSystolicPE_308_io_enable_o;
  wire                uSystolicPE_308_io_clear_o;
  wire                uSystolicPE_309_io_mac_done;
  wire                uSystolicPE_309_io_enable_i;
  wire                uSystolicPE_309_io_clear_i;
  wire                uSystolicPE_309_io_enable_w;
  wire                uSystolicPE_309_io_clear_w;
  wire                uSystolicPE_309_io_enable_o;
  wire                uSystolicPE_309_io_clear_o;
  wire                uSystolicPE_310_io_mac_done;
  wire                uSystolicPE_310_io_enable_i;
  wire                uSystolicPE_310_io_clear_i;
  wire                uSystolicPE_310_io_enable_w;
  wire                uSystolicPE_310_io_clear_w;
  wire                uSystolicPE_310_io_enable_o;
  wire                uSystolicPE_310_io_clear_o;
  wire                uSystolicPE_311_io_mac_done;
  wire                uSystolicPE_311_io_enable_i;
  wire                uSystolicPE_311_io_clear_i;
  wire                uSystolicPE_311_io_enable_w;
  wire                uSystolicPE_311_io_clear_w;
  wire                uSystolicPE_311_io_enable_o;
  wire                uSystolicPE_311_io_clear_o;
  wire                uSystolicPE_312_io_mac_done;
  wire                uSystolicPE_312_io_enable_i;
  wire                uSystolicPE_312_io_clear_i;
  wire                uSystolicPE_312_io_enable_w;
  wire                uSystolicPE_312_io_clear_w;
  wire                uSystolicPE_312_io_enable_o;
  wire                uSystolicPE_312_io_clear_o;
  wire                uSystolicPE_313_io_mac_done;
  wire                uSystolicPE_313_io_enable_i;
  wire                uSystolicPE_313_io_clear_i;
  wire                uSystolicPE_313_io_enable_w;
  wire                uSystolicPE_313_io_clear_w;
  wire                uSystolicPE_313_io_enable_o;
  wire                uSystolicPE_313_io_clear_o;
  wire                uSystolicPE_314_io_mac_done;
  wire                uSystolicPE_314_io_enable_i;
  wire                uSystolicPE_314_io_clear_i;
  wire                uSystolicPE_314_io_enable_w;
  wire                uSystolicPE_314_io_clear_w;
  wire                uSystolicPE_314_io_enable_o;
  wire                uSystolicPE_314_io_clear_o;
  wire                uSystolicPEBorder_21_io_mac_done;
  wire                uSystolicPEBorder_21_io_enable_i;
  wire                uSystolicPEBorder_21_io_clear_i;
  wire                uSystolicPEBorder_21_io_enable_w;
  wire                uSystolicPEBorder_21_io_clear_w;
  wire                uSystolicPEBorder_21_io_enable_o;
  wire                uSystolicPEBorder_21_io_clear_o;
  wire                uSystolicPE_315_io_mac_done;
  wire                uSystolicPE_315_io_enable_i;
  wire                uSystolicPE_315_io_clear_i;
  wire                uSystolicPE_315_io_enable_w;
  wire                uSystolicPE_315_io_clear_w;
  wire                uSystolicPE_315_io_enable_o;
  wire                uSystolicPE_315_io_clear_o;
  wire                uSystolicPE_316_io_mac_done;
  wire                uSystolicPE_316_io_enable_i;
  wire                uSystolicPE_316_io_clear_i;
  wire                uSystolicPE_316_io_enable_w;
  wire                uSystolicPE_316_io_clear_w;
  wire                uSystolicPE_316_io_enable_o;
  wire                uSystolicPE_316_io_clear_o;
  wire                uSystolicPE_317_io_mac_done;
  wire                uSystolicPE_317_io_enable_i;
  wire                uSystolicPE_317_io_clear_i;
  wire                uSystolicPE_317_io_enable_w;
  wire                uSystolicPE_317_io_clear_w;
  wire                uSystolicPE_317_io_enable_o;
  wire                uSystolicPE_317_io_clear_o;
  wire                uSystolicPE_318_io_mac_done;
  wire                uSystolicPE_318_io_enable_i;
  wire                uSystolicPE_318_io_clear_i;
  wire                uSystolicPE_318_io_enable_w;
  wire                uSystolicPE_318_io_clear_w;
  wire                uSystolicPE_318_io_enable_o;
  wire                uSystolicPE_318_io_clear_o;
  wire                uSystolicPE_319_io_mac_done;
  wire                uSystolicPE_319_io_enable_i;
  wire                uSystolicPE_319_io_clear_i;
  wire                uSystolicPE_319_io_enable_w;
  wire                uSystolicPE_319_io_clear_w;
  wire                uSystolicPE_319_io_enable_o;
  wire                uSystolicPE_319_io_clear_o;
  wire                uSystolicPE_320_io_mac_done;
  wire                uSystolicPE_320_io_enable_i;
  wire                uSystolicPE_320_io_clear_i;
  wire                uSystolicPE_320_io_enable_w;
  wire                uSystolicPE_320_io_clear_w;
  wire                uSystolicPE_320_io_enable_o;
  wire                uSystolicPE_320_io_clear_o;
  wire                uSystolicPE_321_io_mac_done;
  wire                uSystolicPE_321_io_enable_i;
  wire                uSystolicPE_321_io_clear_i;
  wire                uSystolicPE_321_io_enable_w;
  wire                uSystolicPE_321_io_clear_w;
  wire                uSystolicPE_321_io_enable_o;
  wire                uSystolicPE_321_io_clear_o;
  wire                uSystolicPE_322_io_mac_done;
  wire                uSystolicPE_322_io_enable_i;
  wire                uSystolicPE_322_io_clear_i;
  wire                uSystolicPE_322_io_enable_w;
  wire                uSystolicPE_322_io_clear_w;
  wire                uSystolicPE_322_io_enable_o;
  wire                uSystolicPE_322_io_clear_o;
  wire                uSystolicPE_323_io_mac_done;
  wire                uSystolicPE_323_io_enable_i;
  wire                uSystolicPE_323_io_clear_i;
  wire                uSystolicPE_323_io_enable_w;
  wire                uSystolicPE_323_io_clear_w;
  wire                uSystolicPE_323_io_enable_o;
  wire                uSystolicPE_323_io_clear_o;
  wire                uSystolicPE_324_io_mac_done;
  wire                uSystolicPE_324_io_enable_i;
  wire                uSystolicPE_324_io_clear_i;
  wire                uSystolicPE_324_io_enable_w;
  wire                uSystolicPE_324_io_clear_w;
  wire                uSystolicPE_324_io_enable_o;
  wire                uSystolicPE_324_io_clear_o;
  wire                uSystolicPE_325_io_mac_done;
  wire                uSystolicPE_325_io_enable_i;
  wire                uSystolicPE_325_io_clear_i;
  wire                uSystolicPE_325_io_enable_w;
  wire                uSystolicPE_325_io_clear_w;
  wire                uSystolicPE_325_io_enable_o;
  wire                uSystolicPE_325_io_clear_o;
  wire                uSystolicPE_326_io_mac_done;
  wire                uSystolicPE_326_io_enable_i;
  wire                uSystolicPE_326_io_clear_i;
  wire                uSystolicPE_326_io_enable_w;
  wire                uSystolicPE_326_io_clear_w;
  wire                uSystolicPE_326_io_enable_o;
  wire                uSystolicPE_326_io_clear_o;
  wire                uSystolicPE_327_io_mac_done;
  wire                uSystolicPE_327_io_enable_i;
  wire                uSystolicPE_327_io_clear_i;
  wire                uSystolicPE_327_io_enable_w;
  wire                uSystolicPE_327_io_clear_w;
  wire                uSystolicPE_327_io_enable_o;
  wire                uSystolicPE_327_io_clear_o;
  wire                uSystolicPE_328_io_mac_done;
  wire                uSystolicPE_328_io_enable_i;
  wire                uSystolicPE_328_io_clear_i;
  wire                uSystolicPE_328_io_enable_w;
  wire                uSystolicPE_328_io_clear_w;
  wire                uSystolicPE_328_io_enable_o;
  wire                uSystolicPE_328_io_clear_o;
  wire                uSystolicPE_329_io_mac_done;
  wire                uSystolicPE_329_io_enable_i;
  wire                uSystolicPE_329_io_clear_i;
  wire                uSystolicPE_329_io_enable_w;
  wire                uSystolicPE_329_io_clear_w;
  wire                uSystolicPE_329_io_enable_o;
  wire                uSystolicPE_329_io_clear_o;
  wire                uSystolicPEBorder_22_io_mac_done;
  wire                uSystolicPEBorder_22_io_enable_i;
  wire                uSystolicPEBorder_22_io_clear_i;
  wire                uSystolicPEBorder_22_io_enable_w;
  wire                uSystolicPEBorder_22_io_clear_w;
  wire                uSystolicPEBorder_22_io_enable_o;
  wire                uSystolicPEBorder_22_io_clear_o;
  wire                uSystolicPE_330_io_mac_done;
  wire                uSystolicPE_330_io_enable_i;
  wire                uSystolicPE_330_io_clear_i;
  wire                uSystolicPE_330_io_enable_w;
  wire                uSystolicPE_330_io_clear_w;
  wire                uSystolicPE_330_io_enable_o;
  wire                uSystolicPE_330_io_clear_o;
  wire                uSystolicPE_331_io_mac_done;
  wire                uSystolicPE_331_io_enable_i;
  wire                uSystolicPE_331_io_clear_i;
  wire                uSystolicPE_331_io_enable_w;
  wire                uSystolicPE_331_io_clear_w;
  wire                uSystolicPE_331_io_enable_o;
  wire                uSystolicPE_331_io_clear_o;
  wire                uSystolicPE_332_io_mac_done;
  wire                uSystolicPE_332_io_enable_i;
  wire                uSystolicPE_332_io_clear_i;
  wire                uSystolicPE_332_io_enable_w;
  wire                uSystolicPE_332_io_clear_w;
  wire                uSystolicPE_332_io_enable_o;
  wire                uSystolicPE_332_io_clear_o;
  wire                uSystolicPE_333_io_mac_done;
  wire                uSystolicPE_333_io_enable_i;
  wire                uSystolicPE_333_io_clear_i;
  wire                uSystolicPE_333_io_enable_w;
  wire                uSystolicPE_333_io_clear_w;
  wire                uSystolicPE_333_io_enable_o;
  wire                uSystolicPE_333_io_clear_o;
  wire                uSystolicPE_334_io_mac_done;
  wire                uSystolicPE_334_io_enable_i;
  wire                uSystolicPE_334_io_clear_i;
  wire                uSystolicPE_334_io_enable_w;
  wire                uSystolicPE_334_io_clear_w;
  wire                uSystolicPE_334_io_enable_o;
  wire                uSystolicPE_334_io_clear_o;
  wire                uSystolicPE_335_io_mac_done;
  wire                uSystolicPE_335_io_enable_i;
  wire                uSystolicPE_335_io_clear_i;
  wire                uSystolicPE_335_io_enable_w;
  wire                uSystolicPE_335_io_clear_w;
  wire                uSystolicPE_335_io_enable_o;
  wire                uSystolicPE_335_io_clear_o;
  wire                uSystolicPE_336_io_mac_done;
  wire                uSystolicPE_336_io_enable_i;
  wire                uSystolicPE_336_io_clear_i;
  wire                uSystolicPE_336_io_enable_w;
  wire                uSystolicPE_336_io_clear_w;
  wire                uSystolicPE_336_io_enable_o;
  wire                uSystolicPE_336_io_clear_o;
  wire                uSystolicPE_337_io_mac_done;
  wire                uSystolicPE_337_io_enable_i;
  wire                uSystolicPE_337_io_clear_i;
  wire                uSystolicPE_337_io_enable_w;
  wire                uSystolicPE_337_io_clear_w;
  wire                uSystolicPE_337_io_enable_o;
  wire                uSystolicPE_337_io_clear_o;
  wire                uSystolicPE_338_io_mac_done;
  wire                uSystolicPE_338_io_enable_i;
  wire                uSystolicPE_338_io_clear_i;
  wire                uSystolicPE_338_io_enable_w;
  wire                uSystolicPE_338_io_clear_w;
  wire                uSystolicPE_338_io_enable_o;
  wire                uSystolicPE_338_io_clear_o;
  wire                uSystolicPE_339_io_mac_done;
  wire                uSystolicPE_339_io_enable_i;
  wire                uSystolicPE_339_io_clear_i;
  wire                uSystolicPE_339_io_enable_w;
  wire                uSystolicPE_339_io_clear_w;
  wire                uSystolicPE_339_io_enable_o;
  wire                uSystolicPE_339_io_clear_o;
  wire                uSystolicPE_340_io_mac_done;
  wire                uSystolicPE_340_io_enable_i;
  wire                uSystolicPE_340_io_clear_i;
  wire                uSystolicPE_340_io_enable_w;
  wire                uSystolicPE_340_io_clear_w;
  wire                uSystolicPE_340_io_enable_o;
  wire                uSystolicPE_340_io_clear_o;
  wire                uSystolicPE_341_io_mac_done;
  wire                uSystolicPE_341_io_enable_i;
  wire                uSystolicPE_341_io_clear_i;
  wire                uSystolicPE_341_io_enable_w;
  wire                uSystolicPE_341_io_clear_w;
  wire                uSystolicPE_341_io_enable_o;
  wire                uSystolicPE_341_io_clear_o;
  wire                uSystolicPE_342_io_mac_done;
  wire                uSystolicPE_342_io_enable_i;
  wire                uSystolicPE_342_io_clear_i;
  wire                uSystolicPE_342_io_enable_w;
  wire                uSystolicPE_342_io_clear_w;
  wire                uSystolicPE_342_io_enable_o;
  wire                uSystolicPE_342_io_clear_o;
  wire                uSystolicPE_343_io_mac_done;
  wire                uSystolicPE_343_io_enable_i;
  wire                uSystolicPE_343_io_clear_i;
  wire                uSystolicPE_343_io_enable_w;
  wire                uSystolicPE_343_io_clear_w;
  wire                uSystolicPE_343_io_enable_o;
  wire                uSystolicPE_343_io_clear_o;
  wire                uSystolicPE_344_io_mac_done;
  wire                uSystolicPE_344_io_enable_i;
  wire                uSystolicPE_344_io_clear_i;
  wire                uSystolicPE_344_io_enable_w;
  wire                uSystolicPE_344_io_clear_w;
  wire                uSystolicPE_344_io_enable_o;
  wire                uSystolicPE_344_io_clear_o;
  wire                uSystolicPEBorder_23_io_mac_done;
  wire                uSystolicPEBorder_23_io_enable_i;
  wire                uSystolicPEBorder_23_io_clear_i;
  wire                uSystolicPEBorder_23_io_enable_w;
  wire                uSystolicPEBorder_23_io_clear_w;
  wire                uSystolicPEBorder_23_io_enable_o;
  wire                uSystolicPEBorder_23_io_clear_o;
  wire                uSystolicPE_345_io_mac_done;
  wire                uSystolicPE_345_io_enable_i;
  wire                uSystolicPE_345_io_clear_i;
  wire                uSystolicPE_345_io_enable_w;
  wire                uSystolicPE_345_io_clear_w;
  wire                uSystolicPE_345_io_enable_o;
  wire                uSystolicPE_345_io_clear_o;
  wire                uSystolicPE_346_io_mac_done;
  wire                uSystolicPE_346_io_enable_i;
  wire                uSystolicPE_346_io_clear_i;
  wire                uSystolicPE_346_io_enable_w;
  wire                uSystolicPE_346_io_clear_w;
  wire                uSystolicPE_346_io_enable_o;
  wire                uSystolicPE_346_io_clear_o;
  wire                uSystolicPE_347_io_mac_done;
  wire                uSystolicPE_347_io_enable_i;
  wire                uSystolicPE_347_io_clear_i;
  wire                uSystolicPE_347_io_enable_w;
  wire                uSystolicPE_347_io_clear_w;
  wire                uSystolicPE_347_io_enable_o;
  wire                uSystolicPE_347_io_clear_o;
  wire                uSystolicPE_348_io_mac_done;
  wire                uSystolicPE_348_io_enable_i;
  wire                uSystolicPE_348_io_clear_i;
  wire                uSystolicPE_348_io_enable_w;
  wire                uSystolicPE_348_io_clear_w;
  wire                uSystolicPE_348_io_enable_o;
  wire                uSystolicPE_348_io_clear_o;
  wire                uSystolicPE_349_io_mac_done;
  wire                uSystolicPE_349_io_enable_i;
  wire                uSystolicPE_349_io_clear_i;
  wire                uSystolicPE_349_io_enable_w;
  wire                uSystolicPE_349_io_clear_w;
  wire                uSystolicPE_349_io_enable_o;
  wire                uSystolicPE_349_io_clear_o;
  wire                uSystolicPE_350_io_mac_done;
  wire                uSystolicPE_350_io_enable_i;
  wire                uSystolicPE_350_io_clear_i;
  wire                uSystolicPE_350_io_enable_w;
  wire                uSystolicPE_350_io_clear_w;
  wire                uSystolicPE_350_io_enable_o;
  wire                uSystolicPE_350_io_clear_o;
  wire                uSystolicPE_351_io_mac_done;
  wire                uSystolicPE_351_io_enable_i;
  wire                uSystolicPE_351_io_clear_i;
  wire                uSystolicPE_351_io_enable_w;
  wire                uSystolicPE_351_io_clear_w;
  wire                uSystolicPE_351_io_enable_o;
  wire                uSystolicPE_351_io_clear_o;
  wire                uSystolicPE_352_io_mac_done;
  wire                uSystolicPE_352_io_enable_i;
  wire                uSystolicPE_352_io_clear_i;
  wire                uSystolicPE_352_io_enable_w;
  wire                uSystolicPE_352_io_clear_w;
  wire                uSystolicPE_352_io_enable_o;
  wire                uSystolicPE_352_io_clear_o;
  wire                uSystolicPE_353_io_mac_done;
  wire                uSystolicPE_353_io_enable_i;
  wire                uSystolicPE_353_io_clear_i;
  wire                uSystolicPE_353_io_enable_w;
  wire                uSystolicPE_353_io_clear_w;
  wire                uSystolicPE_353_io_enable_o;
  wire                uSystolicPE_353_io_clear_o;
  wire                uSystolicPE_354_io_mac_done;
  wire                uSystolicPE_354_io_enable_i;
  wire                uSystolicPE_354_io_clear_i;
  wire                uSystolicPE_354_io_enable_w;
  wire                uSystolicPE_354_io_clear_w;
  wire                uSystolicPE_354_io_enable_o;
  wire                uSystolicPE_354_io_clear_o;
  wire                uSystolicPE_355_io_mac_done;
  wire                uSystolicPE_355_io_enable_i;
  wire                uSystolicPE_355_io_clear_i;
  wire                uSystolicPE_355_io_enable_w;
  wire                uSystolicPE_355_io_clear_w;
  wire                uSystolicPE_355_io_enable_o;
  wire                uSystolicPE_355_io_clear_o;
  wire                uSystolicPE_356_io_mac_done;
  wire                uSystolicPE_356_io_enable_i;
  wire                uSystolicPE_356_io_clear_i;
  wire                uSystolicPE_356_io_enable_w;
  wire                uSystolicPE_356_io_clear_w;
  wire                uSystolicPE_356_io_enable_o;
  wire                uSystolicPE_356_io_clear_o;
  wire                uSystolicPE_357_io_mac_done;
  wire                uSystolicPE_357_io_enable_i;
  wire                uSystolicPE_357_io_clear_i;
  wire                uSystolicPE_357_io_enable_w;
  wire                uSystolicPE_357_io_clear_w;
  wire                uSystolicPE_357_io_enable_o;
  wire                uSystolicPE_357_io_clear_o;
  wire                uSystolicPE_358_io_mac_done;
  wire                uSystolicPE_358_io_enable_i;
  wire                uSystolicPE_358_io_clear_i;
  wire                uSystolicPE_358_io_enable_w;
  wire                uSystolicPE_358_io_clear_w;
  wire                uSystolicPE_358_io_enable_o;
  wire                uSystolicPE_358_io_clear_o;
  wire                uSystolicPE_359_io_mac_done;
  wire                uSystolicPE_359_io_enable_i;
  wire                uSystolicPE_359_io_clear_i;
  wire                uSystolicPE_359_io_enable_w;
  wire                uSystolicPE_359_io_clear_w;
  wire                uSystolicPE_359_io_enable_o;
  wire                uSystolicPE_359_io_clear_o;
  wire                uSystolicPEBorder_24_io_mac_done;
  wire                uSystolicPEBorder_24_io_enable_i;
  wire                uSystolicPEBorder_24_io_clear_i;
  wire                uSystolicPEBorder_24_io_enable_w;
  wire                uSystolicPEBorder_24_io_clear_w;
  wire                uSystolicPEBorder_24_io_enable_o;
  wire                uSystolicPEBorder_24_io_clear_o;
  wire                uSystolicPE_360_io_mac_done;
  wire                uSystolicPE_360_io_enable_i;
  wire                uSystolicPE_360_io_clear_i;
  wire                uSystolicPE_360_io_enable_w;
  wire                uSystolicPE_360_io_clear_w;
  wire                uSystolicPE_360_io_enable_o;
  wire                uSystolicPE_360_io_clear_o;
  wire                uSystolicPE_361_io_mac_done;
  wire                uSystolicPE_361_io_enable_i;
  wire                uSystolicPE_361_io_clear_i;
  wire                uSystolicPE_361_io_enable_w;
  wire                uSystolicPE_361_io_clear_w;
  wire                uSystolicPE_361_io_enable_o;
  wire                uSystolicPE_361_io_clear_o;
  wire                uSystolicPE_362_io_mac_done;
  wire                uSystolicPE_362_io_enable_i;
  wire                uSystolicPE_362_io_clear_i;
  wire                uSystolicPE_362_io_enable_w;
  wire                uSystolicPE_362_io_clear_w;
  wire                uSystolicPE_362_io_enable_o;
  wire                uSystolicPE_362_io_clear_o;
  wire                uSystolicPE_363_io_mac_done;
  wire                uSystolicPE_363_io_enable_i;
  wire                uSystolicPE_363_io_clear_i;
  wire                uSystolicPE_363_io_enable_w;
  wire                uSystolicPE_363_io_clear_w;
  wire                uSystolicPE_363_io_enable_o;
  wire                uSystolicPE_363_io_clear_o;
  wire                uSystolicPE_364_io_mac_done;
  wire                uSystolicPE_364_io_enable_i;
  wire                uSystolicPE_364_io_clear_i;
  wire                uSystolicPE_364_io_enable_w;
  wire                uSystolicPE_364_io_clear_w;
  wire                uSystolicPE_364_io_enable_o;
  wire                uSystolicPE_364_io_clear_o;
  wire                uSystolicPE_365_io_mac_done;
  wire                uSystolicPE_365_io_enable_i;
  wire                uSystolicPE_365_io_clear_i;
  wire                uSystolicPE_365_io_enable_w;
  wire                uSystolicPE_365_io_clear_w;
  wire                uSystolicPE_365_io_enable_o;
  wire                uSystolicPE_365_io_clear_o;
  wire                uSystolicPE_366_io_mac_done;
  wire                uSystolicPE_366_io_enable_i;
  wire                uSystolicPE_366_io_clear_i;
  wire                uSystolicPE_366_io_enable_w;
  wire                uSystolicPE_366_io_clear_w;
  wire                uSystolicPE_366_io_enable_o;
  wire                uSystolicPE_366_io_clear_o;
  wire                uSystolicPE_367_io_mac_done;
  wire                uSystolicPE_367_io_enable_i;
  wire                uSystolicPE_367_io_clear_i;
  wire                uSystolicPE_367_io_enable_w;
  wire                uSystolicPE_367_io_clear_w;
  wire                uSystolicPE_367_io_enable_o;
  wire                uSystolicPE_367_io_clear_o;
  wire                uSystolicPE_368_io_mac_done;
  wire                uSystolicPE_368_io_enable_i;
  wire                uSystolicPE_368_io_clear_i;
  wire                uSystolicPE_368_io_enable_w;
  wire                uSystolicPE_368_io_clear_w;
  wire                uSystolicPE_368_io_enable_o;
  wire                uSystolicPE_368_io_clear_o;
  wire                uSystolicPE_369_io_mac_done;
  wire                uSystolicPE_369_io_enable_i;
  wire                uSystolicPE_369_io_clear_i;
  wire                uSystolicPE_369_io_enable_w;
  wire                uSystolicPE_369_io_clear_w;
  wire                uSystolicPE_369_io_enable_o;
  wire                uSystolicPE_369_io_clear_o;
  wire                uSystolicPE_370_io_mac_done;
  wire                uSystolicPE_370_io_enable_i;
  wire                uSystolicPE_370_io_clear_i;
  wire                uSystolicPE_370_io_enable_w;
  wire                uSystolicPE_370_io_clear_w;
  wire                uSystolicPE_370_io_enable_o;
  wire                uSystolicPE_370_io_clear_o;
  wire                uSystolicPE_371_io_mac_done;
  wire                uSystolicPE_371_io_enable_i;
  wire                uSystolicPE_371_io_clear_i;
  wire                uSystolicPE_371_io_enable_w;
  wire                uSystolicPE_371_io_clear_w;
  wire                uSystolicPE_371_io_enable_o;
  wire                uSystolicPE_371_io_clear_o;
  wire                uSystolicPE_372_io_mac_done;
  wire                uSystolicPE_372_io_enable_i;
  wire                uSystolicPE_372_io_clear_i;
  wire                uSystolicPE_372_io_enable_w;
  wire                uSystolicPE_372_io_clear_w;
  wire                uSystolicPE_372_io_enable_o;
  wire                uSystolicPE_372_io_clear_o;
  wire                uSystolicPE_373_io_mac_done;
  wire                uSystolicPE_373_io_enable_i;
  wire                uSystolicPE_373_io_clear_i;
  wire                uSystolicPE_373_io_enable_w;
  wire                uSystolicPE_373_io_clear_w;
  wire                uSystolicPE_373_io_enable_o;
  wire                uSystolicPE_373_io_clear_o;
  wire                uSystolicPE_374_io_mac_done;
  wire                uSystolicPE_374_io_enable_i;
  wire                uSystolicPE_374_io_clear_i;
  wire                uSystolicPE_374_io_enable_w;
  wire                uSystolicPE_374_io_clear_w;
  wire                uSystolicPE_374_io_enable_o;
  wire                uSystolicPE_374_io_clear_o;
  wire                uSystolicPEBorder_25_io_mac_done;
  wire                uSystolicPEBorder_25_io_enable_i;
  wire                uSystolicPEBorder_25_io_clear_i;
  wire                uSystolicPEBorder_25_io_enable_w;
  wire                uSystolicPEBorder_25_io_clear_w;
  wire                uSystolicPEBorder_25_io_enable_o;
  wire                uSystolicPEBorder_25_io_clear_o;
  wire                uSystolicPE_375_io_mac_done;
  wire                uSystolicPE_375_io_enable_i;
  wire                uSystolicPE_375_io_clear_i;
  wire                uSystolicPE_375_io_enable_w;
  wire                uSystolicPE_375_io_clear_w;
  wire                uSystolicPE_375_io_enable_o;
  wire                uSystolicPE_375_io_clear_o;
  wire                uSystolicPE_376_io_mac_done;
  wire                uSystolicPE_376_io_enable_i;
  wire                uSystolicPE_376_io_clear_i;
  wire                uSystolicPE_376_io_enable_w;
  wire                uSystolicPE_376_io_clear_w;
  wire                uSystolicPE_376_io_enable_o;
  wire                uSystolicPE_376_io_clear_o;
  wire                uSystolicPE_377_io_mac_done;
  wire                uSystolicPE_377_io_enable_i;
  wire                uSystolicPE_377_io_clear_i;
  wire                uSystolicPE_377_io_enable_w;
  wire                uSystolicPE_377_io_clear_w;
  wire                uSystolicPE_377_io_enable_o;
  wire                uSystolicPE_377_io_clear_o;
  wire                uSystolicPE_378_io_mac_done;
  wire                uSystolicPE_378_io_enable_i;
  wire                uSystolicPE_378_io_clear_i;
  wire                uSystolicPE_378_io_enable_w;
  wire                uSystolicPE_378_io_clear_w;
  wire                uSystolicPE_378_io_enable_o;
  wire                uSystolicPE_378_io_clear_o;
  wire                uSystolicPE_379_io_mac_done;
  wire                uSystolicPE_379_io_enable_i;
  wire                uSystolicPE_379_io_clear_i;
  wire                uSystolicPE_379_io_enable_w;
  wire                uSystolicPE_379_io_clear_w;
  wire                uSystolicPE_379_io_enable_o;
  wire                uSystolicPE_379_io_clear_o;
  wire                uSystolicPE_380_io_mac_done;
  wire                uSystolicPE_380_io_enable_i;
  wire                uSystolicPE_380_io_clear_i;
  wire                uSystolicPE_380_io_enable_w;
  wire                uSystolicPE_380_io_clear_w;
  wire                uSystolicPE_380_io_enable_o;
  wire                uSystolicPE_380_io_clear_o;
  wire                uSystolicPE_381_io_mac_done;
  wire                uSystolicPE_381_io_enable_i;
  wire                uSystolicPE_381_io_clear_i;
  wire                uSystolicPE_381_io_enable_w;
  wire                uSystolicPE_381_io_clear_w;
  wire                uSystolicPE_381_io_enable_o;
  wire                uSystolicPE_381_io_clear_o;
  wire                uSystolicPE_382_io_mac_done;
  wire                uSystolicPE_382_io_enable_i;
  wire                uSystolicPE_382_io_clear_i;
  wire                uSystolicPE_382_io_enable_w;
  wire                uSystolicPE_382_io_clear_w;
  wire                uSystolicPE_382_io_enable_o;
  wire                uSystolicPE_382_io_clear_o;
  wire                uSystolicPE_383_io_mac_done;
  wire                uSystolicPE_383_io_enable_i;
  wire                uSystolicPE_383_io_clear_i;
  wire                uSystolicPE_383_io_enable_w;
  wire                uSystolicPE_383_io_clear_w;
  wire                uSystolicPE_383_io_enable_o;
  wire                uSystolicPE_383_io_clear_o;
  wire                uSystolicPE_384_io_mac_done;
  wire                uSystolicPE_384_io_enable_i;
  wire                uSystolicPE_384_io_clear_i;
  wire                uSystolicPE_384_io_enable_w;
  wire                uSystolicPE_384_io_clear_w;
  wire                uSystolicPE_384_io_enable_o;
  wire                uSystolicPE_384_io_clear_o;
  wire                uSystolicPE_385_io_mac_done;
  wire                uSystolicPE_385_io_enable_i;
  wire                uSystolicPE_385_io_clear_i;
  wire                uSystolicPE_385_io_enable_w;
  wire                uSystolicPE_385_io_clear_w;
  wire                uSystolicPE_385_io_enable_o;
  wire                uSystolicPE_385_io_clear_o;
  wire                uSystolicPE_386_io_mac_done;
  wire                uSystolicPE_386_io_enable_i;
  wire                uSystolicPE_386_io_clear_i;
  wire                uSystolicPE_386_io_enable_w;
  wire                uSystolicPE_386_io_clear_w;
  wire                uSystolicPE_386_io_enable_o;
  wire                uSystolicPE_386_io_clear_o;
  wire                uSystolicPE_387_io_mac_done;
  wire                uSystolicPE_387_io_enable_i;
  wire                uSystolicPE_387_io_clear_i;
  wire                uSystolicPE_387_io_enable_w;
  wire                uSystolicPE_387_io_clear_w;
  wire                uSystolicPE_387_io_enable_o;
  wire                uSystolicPE_387_io_clear_o;
  wire                uSystolicPE_388_io_mac_done;
  wire                uSystolicPE_388_io_enable_i;
  wire                uSystolicPE_388_io_clear_i;
  wire                uSystolicPE_388_io_enable_w;
  wire                uSystolicPE_388_io_clear_w;
  wire                uSystolicPE_388_io_enable_o;
  wire                uSystolicPE_388_io_clear_o;
  wire                uSystolicPE_389_io_mac_done;
  wire                uSystolicPE_389_io_enable_i;
  wire                uSystolicPE_389_io_clear_i;
  wire                uSystolicPE_389_io_enable_w;
  wire                uSystolicPE_389_io_clear_w;
  wire                uSystolicPE_389_io_enable_o;
  wire                uSystolicPE_389_io_clear_o;
  wire                uSystolicPEBorder_26_io_mac_done;
  wire                uSystolicPEBorder_26_io_enable_i;
  wire                uSystolicPEBorder_26_io_clear_i;
  wire                uSystolicPEBorder_26_io_enable_w;
  wire                uSystolicPEBorder_26_io_clear_w;
  wire                uSystolicPEBorder_26_io_enable_o;
  wire                uSystolicPEBorder_26_io_clear_o;
  wire                uSystolicPE_390_io_mac_done;
  wire                uSystolicPE_390_io_enable_i;
  wire                uSystolicPE_390_io_clear_i;
  wire                uSystolicPE_390_io_enable_w;
  wire                uSystolicPE_390_io_clear_w;
  wire                uSystolicPE_390_io_enable_o;
  wire                uSystolicPE_390_io_clear_o;
  wire                uSystolicPE_391_io_mac_done;
  wire                uSystolicPE_391_io_enable_i;
  wire                uSystolicPE_391_io_clear_i;
  wire                uSystolicPE_391_io_enable_w;
  wire                uSystolicPE_391_io_clear_w;
  wire                uSystolicPE_391_io_enable_o;
  wire                uSystolicPE_391_io_clear_o;
  wire                uSystolicPE_392_io_mac_done;
  wire                uSystolicPE_392_io_enable_i;
  wire                uSystolicPE_392_io_clear_i;
  wire                uSystolicPE_392_io_enable_w;
  wire                uSystolicPE_392_io_clear_w;
  wire                uSystolicPE_392_io_enable_o;
  wire                uSystolicPE_392_io_clear_o;
  wire                uSystolicPE_393_io_mac_done;
  wire                uSystolicPE_393_io_enable_i;
  wire                uSystolicPE_393_io_clear_i;
  wire                uSystolicPE_393_io_enable_w;
  wire                uSystolicPE_393_io_clear_w;
  wire                uSystolicPE_393_io_enable_o;
  wire                uSystolicPE_393_io_clear_o;
  wire                uSystolicPE_394_io_mac_done;
  wire                uSystolicPE_394_io_enable_i;
  wire                uSystolicPE_394_io_clear_i;
  wire                uSystolicPE_394_io_enable_w;
  wire                uSystolicPE_394_io_clear_w;
  wire                uSystolicPE_394_io_enable_o;
  wire                uSystolicPE_394_io_clear_o;
  wire                uSystolicPE_395_io_mac_done;
  wire                uSystolicPE_395_io_enable_i;
  wire                uSystolicPE_395_io_clear_i;
  wire                uSystolicPE_395_io_enable_w;
  wire                uSystolicPE_395_io_clear_w;
  wire                uSystolicPE_395_io_enable_o;
  wire                uSystolicPE_395_io_clear_o;
  wire                uSystolicPE_396_io_mac_done;
  wire                uSystolicPE_396_io_enable_i;
  wire                uSystolicPE_396_io_clear_i;
  wire                uSystolicPE_396_io_enable_w;
  wire                uSystolicPE_396_io_clear_w;
  wire                uSystolicPE_396_io_enable_o;
  wire                uSystolicPE_396_io_clear_o;
  wire                uSystolicPE_397_io_mac_done;
  wire                uSystolicPE_397_io_enable_i;
  wire                uSystolicPE_397_io_clear_i;
  wire                uSystolicPE_397_io_enable_w;
  wire                uSystolicPE_397_io_clear_w;
  wire                uSystolicPE_397_io_enable_o;
  wire                uSystolicPE_397_io_clear_o;
  wire                uSystolicPE_398_io_mac_done;
  wire                uSystolicPE_398_io_enable_i;
  wire                uSystolicPE_398_io_clear_i;
  wire                uSystolicPE_398_io_enable_w;
  wire                uSystolicPE_398_io_clear_w;
  wire                uSystolicPE_398_io_enable_o;
  wire                uSystolicPE_398_io_clear_o;
  wire                uSystolicPE_399_io_mac_done;
  wire                uSystolicPE_399_io_enable_i;
  wire                uSystolicPE_399_io_clear_i;
  wire                uSystolicPE_399_io_enable_w;
  wire                uSystolicPE_399_io_clear_w;
  wire                uSystolicPE_399_io_enable_o;
  wire                uSystolicPE_399_io_clear_o;
  wire                uSystolicPE_400_io_mac_done;
  wire                uSystolicPE_400_io_enable_i;
  wire                uSystolicPE_400_io_clear_i;
  wire                uSystolicPE_400_io_enable_w;
  wire                uSystolicPE_400_io_clear_w;
  wire                uSystolicPE_400_io_enable_o;
  wire                uSystolicPE_400_io_clear_o;
  wire                uSystolicPE_401_io_mac_done;
  wire                uSystolicPE_401_io_enable_i;
  wire                uSystolicPE_401_io_clear_i;
  wire                uSystolicPE_401_io_enable_w;
  wire                uSystolicPE_401_io_clear_w;
  wire                uSystolicPE_401_io_enable_o;
  wire                uSystolicPE_401_io_clear_o;
  wire                uSystolicPE_402_io_mac_done;
  wire                uSystolicPE_402_io_enable_i;
  wire                uSystolicPE_402_io_clear_i;
  wire                uSystolicPE_402_io_enable_w;
  wire                uSystolicPE_402_io_clear_w;
  wire                uSystolicPE_402_io_enable_o;
  wire                uSystolicPE_402_io_clear_o;
  wire                uSystolicPE_403_io_mac_done;
  wire                uSystolicPE_403_io_enable_i;
  wire                uSystolicPE_403_io_clear_i;
  wire                uSystolicPE_403_io_enable_w;
  wire                uSystolicPE_403_io_clear_w;
  wire                uSystolicPE_403_io_enable_o;
  wire                uSystolicPE_403_io_clear_o;
  wire                uSystolicPE_404_io_mac_done;
  wire                uSystolicPE_404_io_enable_i;
  wire                uSystolicPE_404_io_clear_i;
  wire                uSystolicPE_404_io_enable_w;
  wire                uSystolicPE_404_io_clear_w;
  wire                uSystolicPE_404_io_enable_o;
  wire                uSystolicPE_404_io_clear_o;
  wire                uSystolicPEBorder_27_io_mac_done;
  wire                uSystolicPEBorder_27_io_enable_i;
  wire                uSystolicPEBorder_27_io_clear_i;
  wire                uSystolicPEBorder_27_io_enable_w;
  wire                uSystolicPEBorder_27_io_clear_w;
  wire                uSystolicPEBorder_27_io_enable_o;
  wire                uSystolicPEBorder_27_io_clear_o;
  wire                uSystolicPE_405_io_mac_done;
  wire                uSystolicPE_405_io_enable_i;
  wire                uSystolicPE_405_io_clear_i;
  wire                uSystolicPE_405_io_enable_w;
  wire                uSystolicPE_405_io_clear_w;
  wire                uSystolicPE_405_io_enable_o;
  wire                uSystolicPE_405_io_clear_o;
  wire                uSystolicPE_406_io_mac_done;
  wire                uSystolicPE_406_io_enable_i;
  wire                uSystolicPE_406_io_clear_i;
  wire                uSystolicPE_406_io_enable_w;
  wire                uSystolicPE_406_io_clear_w;
  wire                uSystolicPE_406_io_enable_o;
  wire                uSystolicPE_406_io_clear_o;
  wire                uSystolicPE_407_io_mac_done;
  wire                uSystolicPE_407_io_enable_i;
  wire                uSystolicPE_407_io_clear_i;
  wire                uSystolicPE_407_io_enable_w;
  wire                uSystolicPE_407_io_clear_w;
  wire                uSystolicPE_407_io_enable_o;
  wire                uSystolicPE_407_io_clear_o;
  wire                uSystolicPE_408_io_mac_done;
  wire                uSystolicPE_408_io_enable_i;
  wire                uSystolicPE_408_io_clear_i;
  wire                uSystolicPE_408_io_enable_w;
  wire                uSystolicPE_408_io_clear_w;
  wire                uSystolicPE_408_io_enable_o;
  wire                uSystolicPE_408_io_clear_o;
  wire                uSystolicPE_409_io_mac_done;
  wire                uSystolicPE_409_io_enable_i;
  wire                uSystolicPE_409_io_clear_i;
  wire                uSystolicPE_409_io_enable_w;
  wire                uSystolicPE_409_io_clear_w;
  wire                uSystolicPE_409_io_enable_o;
  wire                uSystolicPE_409_io_clear_o;
  wire                uSystolicPE_410_io_mac_done;
  wire                uSystolicPE_410_io_enable_i;
  wire                uSystolicPE_410_io_clear_i;
  wire                uSystolicPE_410_io_enable_w;
  wire                uSystolicPE_410_io_clear_w;
  wire                uSystolicPE_410_io_enable_o;
  wire                uSystolicPE_410_io_clear_o;
  wire                uSystolicPE_411_io_mac_done;
  wire                uSystolicPE_411_io_enable_i;
  wire                uSystolicPE_411_io_clear_i;
  wire                uSystolicPE_411_io_enable_w;
  wire                uSystolicPE_411_io_clear_w;
  wire                uSystolicPE_411_io_enable_o;
  wire                uSystolicPE_411_io_clear_o;
  wire                uSystolicPE_412_io_mac_done;
  wire                uSystolicPE_412_io_enable_i;
  wire                uSystolicPE_412_io_clear_i;
  wire                uSystolicPE_412_io_enable_w;
  wire                uSystolicPE_412_io_clear_w;
  wire                uSystolicPE_412_io_enable_o;
  wire                uSystolicPE_412_io_clear_o;
  wire                uSystolicPE_413_io_mac_done;
  wire                uSystolicPE_413_io_enable_i;
  wire                uSystolicPE_413_io_clear_i;
  wire                uSystolicPE_413_io_enable_w;
  wire                uSystolicPE_413_io_clear_w;
  wire                uSystolicPE_413_io_enable_o;
  wire                uSystolicPE_413_io_clear_o;
  wire                uSystolicPE_414_io_mac_done;
  wire                uSystolicPE_414_io_enable_i;
  wire                uSystolicPE_414_io_clear_i;
  wire                uSystolicPE_414_io_enable_w;
  wire                uSystolicPE_414_io_clear_w;
  wire                uSystolicPE_414_io_enable_o;
  wire                uSystolicPE_414_io_clear_o;
  wire                uSystolicPE_415_io_mac_done;
  wire                uSystolicPE_415_io_enable_i;
  wire                uSystolicPE_415_io_clear_i;
  wire                uSystolicPE_415_io_enable_w;
  wire                uSystolicPE_415_io_clear_w;
  wire                uSystolicPE_415_io_enable_o;
  wire                uSystolicPE_415_io_clear_o;
  wire                uSystolicPE_416_io_mac_done;
  wire                uSystolicPE_416_io_enable_i;
  wire                uSystolicPE_416_io_clear_i;
  wire                uSystolicPE_416_io_enable_w;
  wire                uSystolicPE_416_io_clear_w;
  wire                uSystolicPE_416_io_enable_o;
  wire                uSystolicPE_416_io_clear_o;
  wire                uSystolicPE_417_io_mac_done;
  wire                uSystolicPE_417_io_enable_i;
  wire                uSystolicPE_417_io_clear_i;
  wire                uSystolicPE_417_io_enable_w;
  wire                uSystolicPE_417_io_clear_w;
  wire                uSystolicPE_417_io_enable_o;
  wire                uSystolicPE_417_io_clear_o;
  wire                uSystolicPE_418_io_mac_done;
  wire                uSystolicPE_418_io_enable_i;
  wire                uSystolicPE_418_io_clear_i;
  wire                uSystolicPE_418_io_enable_w;
  wire                uSystolicPE_418_io_clear_w;
  wire                uSystolicPE_418_io_enable_o;
  wire                uSystolicPE_418_io_clear_o;
  wire                uSystolicPE_419_io_mac_done;
  wire                uSystolicPE_419_io_enable_i;
  wire                uSystolicPE_419_io_clear_i;
  wire                uSystolicPE_419_io_enable_w;
  wire                uSystolicPE_419_io_clear_w;
  wire                uSystolicPE_419_io_enable_o;
  wire                uSystolicPE_419_io_clear_o;
  wire                uSystolicPEBorder_28_io_mac_done;
  wire                uSystolicPEBorder_28_io_enable_i;
  wire                uSystolicPEBorder_28_io_clear_i;
  wire                uSystolicPEBorder_28_io_enable_w;
  wire                uSystolicPEBorder_28_io_clear_w;
  wire                uSystolicPEBorder_28_io_enable_o;
  wire                uSystolicPEBorder_28_io_clear_o;
  wire                uSystolicPE_420_io_mac_done;
  wire                uSystolicPE_420_io_enable_i;
  wire                uSystolicPE_420_io_clear_i;
  wire                uSystolicPE_420_io_enable_w;
  wire                uSystolicPE_420_io_clear_w;
  wire                uSystolicPE_420_io_enable_o;
  wire                uSystolicPE_420_io_clear_o;
  wire                uSystolicPE_421_io_mac_done;
  wire                uSystolicPE_421_io_enable_i;
  wire                uSystolicPE_421_io_clear_i;
  wire                uSystolicPE_421_io_enable_w;
  wire                uSystolicPE_421_io_clear_w;
  wire                uSystolicPE_421_io_enable_o;
  wire                uSystolicPE_421_io_clear_o;
  wire                uSystolicPE_422_io_mac_done;
  wire                uSystolicPE_422_io_enable_i;
  wire                uSystolicPE_422_io_clear_i;
  wire                uSystolicPE_422_io_enable_w;
  wire                uSystolicPE_422_io_clear_w;
  wire                uSystolicPE_422_io_enable_o;
  wire                uSystolicPE_422_io_clear_o;
  wire                uSystolicPE_423_io_mac_done;
  wire                uSystolicPE_423_io_enable_i;
  wire                uSystolicPE_423_io_clear_i;
  wire                uSystolicPE_423_io_enable_w;
  wire                uSystolicPE_423_io_clear_w;
  wire                uSystolicPE_423_io_enable_o;
  wire                uSystolicPE_423_io_clear_o;
  wire                uSystolicPE_424_io_mac_done;
  wire                uSystolicPE_424_io_enable_i;
  wire                uSystolicPE_424_io_clear_i;
  wire                uSystolicPE_424_io_enable_w;
  wire                uSystolicPE_424_io_clear_w;
  wire                uSystolicPE_424_io_enable_o;
  wire                uSystolicPE_424_io_clear_o;
  wire                uSystolicPE_425_io_mac_done;
  wire                uSystolicPE_425_io_enable_i;
  wire                uSystolicPE_425_io_clear_i;
  wire                uSystolicPE_425_io_enable_w;
  wire                uSystolicPE_425_io_clear_w;
  wire                uSystolicPE_425_io_enable_o;
  wire                uSystolicPE_425_io_clear_o;
  wire                uSystolicPE_426_io_mac_done;
  wire                uSystolicPE_426_io_enable_i;
  wire                uSystolicPE_426_io_clear_i;
  wire                uSystolicPE_426_io_enable_w;
  wire                uSystolicPE_426_io_clear_w;
  wire                uSystolicPE_426_io_enable_o;
  wire                uSystolicPE_426_io_clear_o;
  wire                uSystolicPE_427_io_mac_done;
  wire                uSystolicPE_427_io_enable_i;
  wire                uSystolicPE_427_io_clear_i;
  wire                uSystolicPE_427_io_enable_w;
  wire                uSystolicPE_427_io_clear_w;
  wire                uSystolicPE_427_io_enable_o;
  wire                uSystolicPE_427_io_clear_o;
  wire                uSystolicPE_428_io_mac_done;
  wire                uSystolicPE_428_io_enable_i;
  wire                uSystolicPE_428_io_clear_i;
  wire                uSystolicPE_428_io_enable_w;
  wire                uSystolicPE_428_io_clear_w;
  wire                uSystolicPE_428_io_enable_o;
  wire                uSystolicPE_428_io_clear_o;
  wire                uSystolicPE_429_io_mac_done;
  wire                uSystolicPE_429_io_enable_i;
  wire                uSystolicPE_429_io_clear_i;
  wire                uSystolicPE_429_io_enable_w;
  wire                uSystolicPE_429_io_clear_w;
  wire                uSystolicPE_429_io_enable_o;
  wire                uSystolicPE_429_io_clear_o;
  wire                uSystolicPE_430_io_mac_done;
  wire                uSystolicPE_430_io_enable_i;
  wire                uSystolicPE_430_io_clear_i;
  wire                uSystolicPE_430_io_enable_w;
  wire                uSystolicPE_430_io_clear_w;
  wire                uSystolicPE_430_io_enable_o;
  wire                uSystolicPE_430_io_clear_o;
  wire                uSystolicPE_431_io_mac_done;
  wire                uSystolicPE_431_io_enable_i;
  wire                uSystolicPE_431_io_clear_i;
  wire                uSystolicPE_431_io_enable_w;
  wire                uSystolicPE_431_io_clear_w;
  wire                uSystolicPE_431_io_enable_o;
  wire                uSystolicPE_431_io_clear_o;
  wire                uSystolicPE_432_io_mac_done;
  wire                uSystolicPE_432_io_enable_i;
  wire                uSystolicPE_432_io_clear_i;
  wire                uSystolicPE_432_io_enable_w;
  wire                uSystolicPE_432_io_clear_w;
  wire                uSystolicPE_432_io_enable_o;
  wire                uSystolicPE_432_io_clear_o;
  wire                uSystolicPE_433_io_mac_done;
  wire                uSystolicPE_433_io_enable_i;
  wire                uSystolicPE_433_io_clear_i;
  wire                uSystolicPE_433_io_enable_w;
  wire                uSystolicPE_433_io_clear_w;
  wire                uSystolicPE_433_io_enable_o;
  wire                uSystolicPE_433_io_clear_o;
  wire                uSystolicPE_434_io_mac_done;
  wire                uSystolicPE_434_io_enable_i;
  wire                uSystolicPE_434_io_clear_i;
  wire                uSystolicPE_434_io_enable_w;
  wire                uSystolicPE_434_io_clear_w;
  wire                uSystolicPE_434_io_enable_o;
  wire                uSystolicPE_434_io_clear_o;
  wire                uSystolicPEBorder_29_io_mac_done;
  wire                uSystolicPEBorder_29_io_enable_i;
  wire                uSystolicPEBorder_29_io_clear_i;
  wire                uSystolicPEBorder_29_io_enable_w;
  wire                uSystolicPEBorder_29_io_clear_w;
  wire                uSystolicPEBorder_29_io_enable_o;
  wire                uSystolicPEBorder_29_io_clear_o;
  wire                uSystolicPE_435_io_mac_done;
  wire                uSystolicPE_435_io_enable_i;
  wire                uSystolicPE_435_io_clear_i;
  wire                uSystolicPE_435_io_enable_w;
  wire                uSystolicPE_435_io_clear_w;
  wire                uSystolicPE_435_io_enable_o;
  wire                uSystolicPE_435_io_clear_o;
  wire                uSystolicPE_436_io_mac_done;
  wire                uSystolicPE_436_io_enable_i;
  wire                uSystolicPE_436_io_clear_i;
  wire                uSystolicPE_436_io_enable_w;
  wire                uSystolicPE_436_io_clear_w;
  wire                uSystolicPE_436_io_enable_o;
  wire                uSystolicPE_436_io_clear_o;
  wire                uSystolicPE_437_io_mac_done;
  wire                uSystolicPE_437_io_enable_i;
  wire                uSystolicPE_437_io_clear_i;
  wire                uSystolicPE_437_io_enable_w;
  wire                uSystolicPE_437_io_clear_w;
  wire                uSystolicPE_437_io_enable_o;
  wire                uSystolicPE_437_io_clear_o;
  wire                uSystolicPE_438_io_mac_done;
  wire                uSystolicPE_438_io_enable_i;
  wire                uSystolicPE_438_io_clear_i;
  wire                uSystolicPE_438_io_enable_w;
  wire                uSystolicPE_438_io_clear_w;
  wire                uSystolicPE_438_io_enable_o;
  wire                uSystolicPE_438_io_clear_o;
  wire                uSystolicPE_439_io_mac_done;
  wire                uSystolicPE_439_io_enable_i;
  wire                uSystolicPE_439_io_clear_i;
  wire                uSystolicPE_439_io_enable_w;
  wire                uSystolicPE_439_io_clear_w;
  wire                uSystolicPE_439_io_enable_o;
  wire                uSystolicPE_439_io_clear_o;
  wire                uSystolicPE_440_io_mac_done;
  wire                uSystolicPE_440_io_enable_i;
  wire                uSystolicPE_440_io_clear_i;
  wire                uSystolicPE_440_io_enable_w;
  wire                uSystolicPE_440_io_clear_w;
  wire                uSystolicPE_440_io_enable_o;
  wire                uSystolicPE_440_io_clear_o;
  wire                uSystolicPE_441_io_mac_done;
  wire                uSystolicPE_441_io_enable_i;
  wire                uSystolicPE_441_io_clear_i;
  wire                uSystolicPE_441_io_enable_w;
  wire                uSystolicPE_441_io_clear_w;
  wire                uSystolicPE_441_io_enable_o;
  wire                uSystolicPE_441_io_clear_o;
  wire                uSystolicPE_442_io_mac_done;
  wire                uSystolicPE_442_io_enable_i;
  wire                uSystolicPE_442_io_clear_i;
  wire                uSystolicPE_442_io_enable_w;
  wire                uSystolicPE_442_io_clear_w;
  wire                uSystolicPE_442_io_enable_o;
  wire                uSystolicPE_442_io_clear_o;
  wire                uSystolicPE_443_io_mac_done;
  wire                uSystolicPE_443_io_enable_i;
  wire                uSystolicPE_443_io_clear_i;
  wire                uSystolicPE_443_io_enable_w;
  wire                uSystolicPE_443_io_clear_w;
  wire                uSystolicPE_443_io_enable_o;
  wire                uSystolicPE_443_io_clear_o;
  wire                uSystolicPE_444_io_mac_done;
  wire                uSystolicPE_444_io_enable_i;
  wire                uSystolicPE_444_io_clear_i;
  wire                uSystolicPE_444_io_enable_w;
  wire                uSystolicPE_444_io_clear_w;
  wire                uSystolicPE_444_io_enable_o;
  wire                uSystolicPE_444_io_clear_o;
  wire                uSystolicPE_445_io_mac_done;
  wire                uSystolicPE_445_io_enable_i;
  wire                uSystolicPE_445_io_clear_i;
  wire                uSystolicPE_445_io_enable_w;
  wire                uSystolicPE_445_io_clear_w;
  wire                uSystolicPE_445_io_enable_o;
  wire                uSystolicPE_445_io_clear_o;
  wire                uSystolicPE_446_io_mac_done;
  wire                uSystolicPE_446_io_enable_i;
  wire                uSystolicPE_446_io_clear_i;
  wire                uSystolicPE_446_io_enable_w;
  wire                uSystolicPE_446_io_clear_w;
  wire                uSystolicPE_446_io_enable_o;
  wire                uSystolicPE_446_io_clear_o;
  wire                uSystolicPE_447_io_mac_done;
  wire                uSystolicPE_447_io_enable_i;
  wire                uSystolicPE_447_io_clear_i;
  wire                uSystolicPE_447_io_enable_w;
  wire                uSystolicPE_447_io_clear_w;
  wire                uSystolicPE_447_io_enable_o;
  wire                uSystolicPE_447_io_clear_o;
  wire                uSystolicPE_448_io_mac_done;
  wire                uSystolicPE_448_io_enable_i;
  wire                uSystolicPE_448_io_clear_i;
  wire                uSystolicPE_448_io_enable_w;
  wire                uSystolicPE_448_io_clear_w;
  wire                uSystolicPE_448_io_enable_o;
  wire                uSystolicPE_448_io_clear_o;
  wire                uSystolicPE_449_io_mac_done;
  wire                uSystolicPE_449_io_enable_i;
  wire                uSystolicPE_449_io_clear_i;
  wire                uSystolicPE_449_io_enable_w;
  wire                uSystolicPE_449_io_clear_w;
  wire                uSystolicPE_449_io_enable_o;
  wire                uSystolicPE_449_io_clear_o;
  wire                uSystolicPEBorder_30_io_mac_done;
  wire                uSystolicPEBorder_30_io_enable_i;
  wire                uSystolicPEBorder_30_io_clear_i;
  wire                uSystolicPEBorder_30_io_enable_w;
  wire                uSystolicPEBorder_30_io_clear_w;
  wire                uSystolicPEBorder_30_io_enable_o;
  wire                uSystolicPEBorder_30_io_clear_o;
  wire                uSystolicPE_450_io_mac_done;
  wire                uSystolicPE_450_io_enable_i;
  wire                uSystolicPE_450_io_clear_i;
  wire                uSystolicPE_450_io_enable_w;
  wire                uSystolicPE_450_io_clear_w;
  wire                uSystolicPE_450_io_enable_o;
  wire                uSystolicPE_450_io_clear_o;
  wire                uSystolicPE_451_io_mac_done;
  wire                uSystolicPE_451_io_enable_i;
  wire                uSystolicPE_451_io_clear_i;
  wire                uSystolicPE_451_io_enable_w;
  wire                uSystolicPE_451_io_clear_w;
  wire                uSystolicPE_451_io_enable_o;
  wire                uSystolicPE_451_io_clear_o;
  wire                uSystolicPE_452_io_mac_done;
  wire                uSystolicPE_452_io_enable_i;
  wire                uSystolicPE_452_io_clear_i;
  wire                uSystolicPE_452_io_enable_w;
  wire                uSystolicPE_452_io_clear_w;
  wire                uSystolicPE_452_io_enable_o;
  wire                uSystolicPE_452_io_clear_o;
  wire                uSystolicPE_453_io_mac_done;
  wire                uSystolicPE_453_io_enable_i;
  wire                uSystolicPE_453_io_clear_i;
  wire                uSystolicPE_453_io_enable_w;
  wire                uSystolicPE_453_io_clear_w;
  wire                uSystolicPE_453_io_enable_o;
  wire                uSystolicPE_453_io_clear_o;
  wire                uSystolicPE_454_io_mac_done;
  wire                uSystolicPE_454_io_enable_i;
  wire                uSystolicPE_454_io_clear_i;
  wire                uSystolicPE_454_io_enable_w;
  wire                uSystolicPE_454_io_clear_w;
  wire                uSystolicPE_454_io_enable_o;
  wire                uSystolicPE_454_io_clear_o;
  wire                uSystolicPE_455_io_mac_done;
  wire                uSystolicPE_455_io_enable_i;
  wire                uSystolicPE_455_io_clear_i;
  wire                uSystolicPE_455_io_enable_w;
  wire                uSystolicPE_455_io_clear_w;
  wire                uSystolicPE_455_io_enable_o;
  wire                uSystolicPE_455_io_clear_o;
  wire                uSystolicPE_456_io_mac_done;
  wire                uSystolicPE_456_io_enable_i;
  wire                uSystolicPE_456_io_clear_i;
  wire                uSystolicPE_456_io_enable_w;
  wire                uSystolicPE_456_io_clear_w;
  wire                uSystolicPE_456_io_enable_o;
  wire                uSystolicPE_456_io_clear_o;
  wire                uSystolicPE_457_io_mac_done;
  wire                uSystolicPE_457_io_enable_i;
  wire                uSystolicPE_457_io_clear_i;
  wire                uSystolicPE_457_io_enable_w;
  wire                uSystolicPE_457_io_clear_w;
  wire                uSystolicPE_457_io_enable_o;
  wire                uSystolicPE_457_io_clear_o;
  wire                uSystolicPE_458_io_mac_done;
  wire                uSystolicPE_458_io_enable_i;
  wire                uSystolicPE_458_io_clear_i;
  wire                uSystolicPE_458_io_enable_w;
  wire                uSystolicPE_458_io_clear_w;
  wire                uSystolicPE_458_io_enable_o;
  wire                uSystolicPE_458_io_clear_o;
  wire                uSystolicPE_459_io_mac_done;
  wire                uSystolicPE_459_io_enable_i;
  wire                uSystolicPE_459_io_clear_i;
  wire                uSystolicPE_459_io_enable_w;
  wire                uSystolicPE_459_io_clear_w;
  wire                uSystolicPE_459_io_enable_o;
  wire                uSystolicPE_459_io_clear_o;
  wire                uSystolicPE_460_io_mac_done;
  wire                uSystolicPE_460_io_enable_i;
  wire                uSystolicPE_460_io_clear_i;
  wire                uSystolicPE_460_io_enable_w;
  wire                uSystolicPE_460_io_clear_w;
  wire                uSystolicPE_460_io_enable_o;
  wire                uSystolicPE_460_io_clear_o;
  wire                uSystolicPE_461_io_mac_done;
  wire                uSystolicPE_461_io_enable_i;
  wire                uSystolicPE_461_io_clear_i;
  wire                uSystolicPE_461_io_enable_w;
  wire                uSystolicPE_461_io_clear_w;
  wire                uSystolicPE_461_io_enable_o;
  wire                uSystolicPE_461_io_clear_o;
  wire                uSystolicPE_462_io_mac_done;
  wire                uSystolicPE_462_io_enable_i;
  wire                uSystolicPE_462_io_clear_i;
  wire                uSystolicPE_462_io_enable_w;
  wire                uSystolicPE_462_io_clear_w;
  wire                uSystolicPE_462_io_enable_o;
  wire                uSystolicPE_462_io_clear_o;
  wire                uSystolicPE_463_io_mac_done;
  wire                uSystolicPE_463_io_enable_i;
  wire                uSystolicPE_463_io_clear_i;
  wire                uSystolicPE_463_io_enable_w;
  wire                uSystolicPE_463_io_clear_w;
  wire                uSystolicPE_463_io_enable_o;
  wire                uSystolicPE_463_io_clear_o;
  wire                uSystolicPE_464_io_mac_done;
  wire                uSystolicPE_464_io_enable_i;
  wire                uSystolicPE_464_io_clear_i;
  wire                uSystolicPE_464_io_enable_w;
  wire                uSystolicPE_464_io_clear_w;
  wire                uSystolicPE_464_io_enable_o;
  wire                uSystolicPE_464_io_clear_o;
  wire                uSystolicPEBorder_31_io_mac_done;
  wire                uSystolicPEBorder_31_io_enable_i;
  wire                uSystolicPEBorder_31_io_clear_i;
  wire                uSystolicPEBorder_31_io_enable_w;
  wire                uSystolicPEBorder_31_io_clear_w;
  wire                uSystolicPEBorder_31_io_enable_o;
  wire                uSystolicPEBorder_31_io_clear_o;
  wire                uSystolicPE_465_io_mac_done;
  wire                uSystolicPE_465_io_enable_i;
  wire                uSystolicPE_465_io_clear_i;
  wire                uSystolicPE_465_io_enable_w;
  wire                uSystolicPE_465_io_clear_w;
  wire                uSystolicPE_465_io_enable_o;
  wire                uSystolicPE_465_io_clear_o;
  wire                uSystolicPE_466_io_mac_done;
  wire                uSystolicPE_466_io_enable_i;
  wire                uSystolicPE_466_io_clear_i;
  wire                uSystolicPE_466_io_enable_w;
  wire                uSystolicPE_466_io_clear_w;
  wire                uSystolicPE_466_io_enable_o;
  wire                uSystolicPE_466_io_clear_o;
  wire                uSystolicPE_467_io_mac_done;
  wire                uSystolicPE_467_io_enable_i;
  wire                uSystolicPE_467_io_clear_i;
  wire                uSystolicPE_467_io_enable_w;
  wire                uSystolicPE_467_io_clear_w;
  wire                uSystolicPE_467_io_enable_o;
  wire                uSystolicPE_467_io_clear_o;
  wire                uSystolicPE_468_io_mac_done;
  wire                uSystolicPE_468_io_enable_i;
  wire                uSystolicPE_468_io_clear_i;
  wire                uSystolicPE_468_io_enable_w;
  wire                uSystolicPE_468_io_clear_w;
  wire                uSystolicPE_468_io_enable_o;
  wire                uSystolicPE_468_io_clear_o;
  wire                uSystolicPE_469_io_mac_done;
  wire                uSystolicPE_469_io_enable_i;
  wire                uSystolicPE_469_io_clear_i;
  wire                uSystolicPE_469_io_enable_w;
  wire                uSystolicPE_469_io_clear_w;
  wire                uSystolicPE_469_io_enable_o;
  wire                uSystolicPE_469_io_clear_o;
  wire                uSystolicPE_470_io_mac_done;
  wire                uSystolicPE_470_io_enable_i;
  wire                uSystolicPE_470_io_clear_i;
  wire                uSystolicPE_470_io_enable_w;
  wire                uSystolicPE_470_io_clear_w;
  wire                uSystolicPE_470_io_enable_o;
  wire                uSystolicPE_470_io_clear_o;
  wire                uSystolicPE_471_io_mac_done;
  wire                uSystolicPE_471_io_enable_i;
  wire                uSystolicPE_471_io_clear_i;
  wire                uSystolicPE_471_io_enable_w;
  wire                uSystolicPE_471_io_clear_w;
  wire                uSystolicPE_471_io_enable_o;
  wire                uSystolicPE_471_io_clear_o;
  wire                uSystolicPE_472_io_mac_done;
  wire                uSystolicPE_472_io_enable_i;
  wire                uSystolicPE_472_io_clear_i;
  wire                uSystolicPE_472_io_enable_w;
  wire                uSystolicPE_472_io_clear_w;
  wire                uSystolicPE_472_io_enable_o;
  wire                uSystolicPE_472_io_clear_o;
  wire                uSystolicPE_473_io_mac_done;
  wire                uSystolicPE_473_io_enable_i;
  wire                uSystolicPE_473_io_clear_i;
  wire                uSystolicPE_473_io_enable_w;
  wire                uSystolicPE_473_io_clear_w;
  wire                uSystolicPE_473_io_enable_o;
  wire                uSystolicPE_473_io_clear_o;
  wire                uSystolicPE_474_io_mac_done;
  wire                uSystolicPE_474_io_enable_i;
  wire                uSystolicPE_474_io_clear_i;
  wire                uSystolicPE_474_io_enable_w;
  wire                uSystolicPE_474_io_clear_w;
  wire                uSystolicPE_474_io_enable_o;
  wire                uSystolicPE_474_io_clear_o;
  wire                uSystolicPE_475_io_mac_done;
  wire                uSystolicPE_475_io_enable_i;
  wire                uSystolicPE_475_io_clear_i;
  wire                uSystolicPE_475_io_enable_w;
  wire                uSystolicPE_475_io_clear_w;
  wire                uSystolicPE_475_io_enable_o;
  wire                uSystolicPE_475_io_clear_o;
  wire                uSystolicPE_476_io_mac_done;
  wire                uSystolicPE_476_io_enable_i;
  wire                uSystolicPE_476_io_clear_i;
  wire                uSystolicPE_476_io_enable_w;
  wire                uSystolicPE_476_io_clear_w;
  wire                uSystolicPE_476_io_enable_o;
  wire                uSystolicPE_476_io_clear_o;
  wire                uSystolicPE_477_io_mac_done;
  wire                uSystolicPE_477_io_enable_i;
  wire                uSystolicPE_477_io_clear_i;
  wire                uSystolicPE_477_io_enable_w;
  wire                uSystolicPE_477_io_clear_w;
  wire                uSystolicPE_477_io_enable_o;
  wire                uSystolicPE_477_io_clear_o;
  wire                uSystolicPE_478_io_mac_done;
  wire                uSystolicPE_478_io_enable_i;
  wire                uSystolicPE_478_io_clear_i;
  wire                uSystolicPE_478_io_enable_w;
  wire                uSystolicPE_478_io_clear_w;
  wire                uSystolicPE_478_io_enable_o;
  wire                uSystolicPE_478_io_clear_o;
  wire                uSystolicPE_479_io_mac_done;
  wire                uSystolicPE_479_io_enable_i;
  wire                uSystolicPE_479_io_clear_i;
  wire                uSystolicPE_479_io_enable_w;
  wire                uSystolicPE_479_io_clear_w;
  wire                uSystolicPE_479_io_enable_o;
  wire                uSystolicPE_479_io_clear_o;
  wire                uSystolicPEBorder_16_io_mac_done_d;
  wire                uSystolicPEBorder_16_io_enable_i_d;
  wire                uSystolicPEBorder_16_io_clear_i_d;
  wire                uSystolicPEBorder_16_io_enable_w_d;
  wire                uSystolicPEBorder_16_io_clear_w_d;
  wire                uSystolicPEBorder_16_io_enable_o_d;
  wire                uSystolicPEBorder_16_io_clear_o_d;
  wire                uSystolicPEBorder_16_io_ifm_sign_d;
  wire                uSystolicPEBorder_16_io_ifm_dff_d;
  wire                uSystolicPEBorder_16_io_wght_sign_d;
  wire       [14:0]   uSystolicPEBorder_16_io_randW_d;
  wire       [14:0]   uSystolicPEBorder_16_io_wght_abs_d;
  wire       [31:0]   uSystolicPEBorder_16_io_ofm_d;
  wire                uSystolicPE_240_io_mac_done_d;
  wire                uSystolicPE_240_io_enable_i_d;
  wire                uSystolicPE_240_io_clear_i_d;
  wire                uSystolicPE_240_io_enable_w_d;
  wire                uSystolicPE_240_io_clear_w_d;
  wire                uSystolicPE_240_io_enable_o_d;
  wire                uSystolicPE_240_io_clear_o_d;
  wire                uSystolicPE_240_io_ifm_sign_d;
  wire                uSystolicPE_240_io_ifm_dff_d;
  wire                uSystolicPE_240_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_240_io_randW_d;
  wire       [14:0]   uSystolicPE_240_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_240_io_ofm_d;
  wire                uSystolicPE_241_io_mac_done_d;
  wire                uSystolicPE_241_io_enable_i_d;
  wire                uSystolicPE_241_io_clear_i_d;
  wire                uSystolicPE_241_io_enable_w_d;
  wire                uSystolicPE_241_io_clear_w_d;
  wire                uSystolicPE_241_io_enable_o_d;
  wire                uSystolicPE_241_io_clear_o_d;
  wire                uSystolicPE_241_io_ifm_sign_d;
  wire                uSystolicPE_241_io_ifm_dff_d;
  wire                uSystolicPE_241_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_241_io_randW_d;
  wire       [14:0]   uSystolicPE_241_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_241_io_ofm_d;
  wire                uSystolicPE_242_io_mac_done_d;
  wire                uSystolicPE_242_io_enable_i_d;
  wire                uSystolicPE_242_io_clear_i_d;
  wire                uSystolicPE_242_io_enable_w_d;
  wire                uSystolicPE_242_io_clear_w_d;
  wire                uSystolicPE_242_io_enable_o_d;
  wire                uSystolicPE_242_io_clear_o_d;
  wire                uSystolicPE_242_io_ifm_sign_d;
  wire                uSystolicPE_242_io_ifm_dff_d;
  wire                uSystolicPE_242_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_242_io_randW_d;
  wire       [14:0]   uSystolicPE_242_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_242_io_ofm_d;
  wire                uSystolicPE_243_io_mac_done_d;
  wire                uSystolicPE_243_io_enable_i_d;
  wire                uSystolicPE_243_io_clear_i_d;
  wire                uSystolicPE_243_io_enable_w_d;
  wire                uSystolicPE_243_io_clear_w_d;
  wire                uSystolicPE_243_io_enable_o_d;
  wire                uSystolicPE_243_io_clear_o_d;
  wire                uSystolicPE_243_io_ifm_sign_d;
  wire                uSystolicPE_243_io_ifm_dff_d;
  wire                uSystolicPE_243_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_243_io_randW_d;
  wire       [14:0]   uSystolicPE_243_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_243_io_ofm_d;
  wire                uSystolicPE_244_io_mac_done_d;
  wire                uSystolicPE_244_io_enable_i_d;
  wire                uSystolicPE_244_io_clear_i_d;
  wire                uSystolicPE_244_io_enable_w_d;
  wire                uSystolicPE_244_io_clear_w_d;
  wire                uSystolicPE_244_io_enable_o_d;
  wire                uSystolicPE_244_io_clear_o_d;
  wire                uSystolicPE_244_io_ifm_sign_d;
  wire                uSystolicPE_244_io_ifm_dff_d;
  wire                uSystolicPE_244_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_244_io_randW_d;
  wire       [14:0]   uSystolicPE_244_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_244_io_ofm_d;
  wire                uSystolicPE_245_io_mac_done_d;
  wire                uSystolicPE_245_io_enable_i_d;
  wire                uSystolicPE_245_io_clear_i_d;
  wire                uSystolicPE_245_io_enable_w_d;
  wire                uSystolicPE_245_io_clear_w_d;
  wire                uSystolicPE_245_io_enable_o_d;
  wire                uSystolicPE_245_io_clear_o_d;
  wire                uSystolicPE_245_io_ifm_sign_d;
  wire                uSystolicPE_245_io_ifm_dff_d;
  wire                uSystolicPE_245_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_245_io_randW_d;
  wire       [14:0]   uSystolicPE_245_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_245_io_ofm_d;
  wire                uSystolicPE_246_io_mac_done_d;
  wire                uSystolicPE_246_io_enable_i_d;
  wire                uSystolicPE_246_io_clear_i_d;
  wire                uSystolicPE_246_io_enable_w_d;
  wire                uSystolicPE_246_io_clear_w_d;
  wire                uSystolicPE_246_io_enable_o_d;
  wire                uSystolicPE_246_io_clear_o_d;
  wire                uSystolicPE_246_io_ifm_sign_d;
  wire                uSystolicPE_246_io_ifm_dff_d;
  wire                uSystolicPE_246_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_246_io_randW_d;
  wire       [14:0]   uSystolicPE_246_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_246_io_ofm_d;
  wire                uSystolicPE_247_io_mac_done_d;
  wire                uSystolicPE_247_io_enable_i_d;
  wire                uSystolicPE_247_io_clear_i_d;
  wire                uSystolicPE_247_io_enable_w_d;
  wire                uSystolicPE_247_io_clear_w_d;
  wire                uSystolicPE_247_io_enable_o_d;
  wire                uSystolicPE_247_io_clear_o_d;
  wire                uSystolicPE_247_io_ifm_sign_d;
  wire                uSystolicPE_247_io_ifm_dff_d;
  wire                uSystolicPE_247_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_247_io_randW_d;
  wire       [14:0]   uSystolicPE_247_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_247_io_ofm_d;
  wire                uSystolicPE_248_io_mac_done_d;
  wire                uSystolicPE_248_io_enable_i_d;
  wire                uSystolicPE_248_io_clear_i_d;
  wire                uSystolicPE_248_io_enable_w_d;
  wire                uSystolicPE_248_io_clear_w_d;
  wire                uSystolicPE_248_io_enable_o_d;
  wire                uSystolicPE_248_io_clear_o_d;
  wire                uSystolicPE_248_io_ifm_sign_d;
  wire                uSystolicPE_248_io_ifm_dff_d;
  wire                uSystolicPE_248_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_248_io_randW_d;
  wire       [14:0]   uSystolicPE_248_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_248_io_ofm_d;
  wire                uSystolicPE_249_io_mac_done_d;
  wire                uSystolicPE_249_io_enable_i_d;
  wire                uSystolicPE_249_io_clear_i_d;
  wire                uSystolicPE_249_io_enable_w_d;
  wire                uSystolicPE_249_io_clear_w_d;
  wire                uSystolicPE_249_io_enable_o_d;
  wire                uSystolicPE_249_io_clear_o_d;
  wire                uSystolicPE_249_io_ifm_sign_d;
  wire                uSystolicPE_249_io_ifm_dff_d;
  wire                uSystolicPE_249_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_249_io_randW_d;
  wire       [14:0]   uSystolicPE_249_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_249_io_ofm_d;
  wire                uSystolicPE_250_io_mac_done_d;
  wire                uSystolicPE_250_io_enable_i_d;
  wire                uSystolicPE_250_io_clear_i_d;
  wire                uSystolicPE_250_io_enable_w_d;
  wire                uSystolicPE_250_io_clear_w_d;
  wire                uSystolicPE_250_io_enable_o_d;
  wire                uSystolicPE_250_io_clear_o_d;
  wire                uSystolicPE_250_io_ifm_sign_d;
  wire                uSystolicPE_250_io_ifm_dff_d;
  wire                uSystolicPE_250_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_250_io_randW_d;
  wire       [14:0]   uSystolicPE_250_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_250_io_ofm_d;
  wire                uSystolicPE_251_io_mac_done_d;
  wire                uSystolicPE_251_io_enable_i_d;
  wire                uSystolicPE_251_io_clear_i_d;
  wire                uSystolicPE_251_io_enable_w_d;
  wire                uSystolicPE_251_io_clear_w_d;
  wire                uSystolicPE_251_io_enable_o_d;
  wire                uSystolicPE_251_io_clear_o_d;
  wire                uSystolicPE_251_io_ifm_sign_d;
  wire                uSystolicPE_251_io_ifm_dff_d;
  wire                uSystolicPE_251_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_251_io_randW_d;
  wire       [14:0]   uSystolicPE_251_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_251_io_ofm_d;
  wire                uSystolicPE_252_io_mac_done_d;
  wire                uSystolicPE_252_io_enable_i_d;
  wire                uSystolicPE_252_io_clear_i_d;
  wire                uSystolicPE_252_io_enable_w_d;
  wire                uSystolicPE_252_io_clear_w_d;
  wire                uSystolicPE_252_io_enable_o_d;
  wire                uSystolicPE_252_io_clear_o_d;
  wire                uSystolicPE_252_io_ifm_sign_d;
  wire                uSystolicPE_252_io_ifm_dff_d;
  wire                uSystolicPE_252_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_252_io_randW_d;
  wire       [14:0]   uSystolicPE_252_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_252_io_ofm_d;
  wire                uSystolicPE_253_io_mac_done_d;
  wire                uSystolicPE_253_io_enable_i_d;
  wire                uSystolicPE_253_io_clear_i_d;
  wire                uSystolicPE_253_io_enable_w_d;
  wire                uSystolicPE_253_io_clear_w_d;
  wire                uSystolicPE_253_io_enable_o_d;
  wire                uSystolicPE_253_io_clear_o_d;
  wire                uSystolicPE_253_io_ifm_sign_d;
  wire                uSystolicPE_253_io_ifm_dff_d;
  wire                uSystolicPE_253_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_253_io_randW_d;
  wire       [14:0]   uSystolicPE_253_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_253_io_ofm_d;
  wire                uSystolicPE_254_io_mac_done_d;
  wire                uSystolicPE_254_io_enable_i_d;
  wire                uSystolicPE_254_io_clear_i_d;
  wire                uSystolicPE_254_io_enable_w_d;
  wire                uSystolicPE_254_io_clear_w_d;
  wire                uSystolicPE_254_io_enable_o_d;
  wire                uSystolicPE_254_io_clear_o_d;
  wire                uSystolicPE_254_io_ifm_sign_d;
  wire                uSystolicPE_254_io_ifm_dff_d;
  wire                uSystolicPE_254_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_254_io_randW_d;
  wire       [14:0]   uSystolicPE_254_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_254_io_ofm_d;
  wire                uSystolicPEBorder_17_io_mac_done_d;
  wire                uSystolicPEBorder_17_io_enable_i_d;
  wire                uSystolicPEBorder_17_io_clear_i_d;
  wire                uSystolicPEBorder_17_io_enable_w_d;
  wire                uSystolicPEBorder_17_io_clear_w_d;
  wire                uSystolicPEBorder_17_io_enable_o_d;
  wire                uSystolicPEBorder_17_io_clear_o_d;
  wire                uSystolicPEBorder_17_io_ifm_sign_d;
  wire                uSystolicPEBorder_17_io_ifm_dff_d;
  wire                uSystolicPEBorder_17_io_wght_sign_d;
  wire       [14:0]   uSystolicPEBorder_17_io_randW_d;
  wire       [14:0]   uSystolicPEBorder_17_io_wght_abs_d;
  wire       [31:0]   uSystolicPEBorder_17_io_ofm_d;
  wire                uSystolicPE_255_io_mac_done_d;
  wire                uSystolicPE_255_io_enable_i_d;
  wire                uSystolicPE_255_io_clear_i_d;
  wire                uSystolicPE_255_io_enable_w_d;
  wire                uSystolicPE_255_io_clear_w_d;
  wire                uSystolicPE_255_io_enable_o_d;
  wire                uSystolicPE_255_io_clear_o_d;
  wire                uSystolicPE_255_io_ifm_sign_d;
  wire                uSystolicPE_255_io_ifm_dff_d;
  wire                uSystolicPE_255_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_255_io_randW_d;
  wire       [14:0]   uSystolicPE_255_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_255_io_ofm_d;
  wire                uSystolicPE_256_io_mac_done_d;
  wire                uSystolicPE_256_io_enable_i_d;
  wire                uSystolicPE_256_io_clear_i_d;
  wire                uSystolicPE_256_io_enable_w_d;
  wire                uSystolicPE_256_io_clear_w_d;
  wire                uSystolicPE_256_io_enable_o_d;
  wire                uSystolicPE_256_io_clear_o_d;
  wire                uSystolicPE_256_io_ifm_sign_d;
  wire                uSystolicPE_256_io_ifm_dff_d;
  wire                uSystolicPE_256_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_256_io_randW_d;
  wire       [14:0]   uSystolicPE_256_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_256_io_ofm_d;
  wire                uSystolicPE_257_io_mac_done_d;
  wire                uSystolicPE_257_io_enable_i_d;
  wire                uSystolicPE_257_io_clear_i_d;
  wire                uSystolicPE_257_io_enable_w_d;
  wire                uSystolicPE_257_io_clear_w_d;
  wire                uSystolicPE_257_io_enable_o_d;
  wire                uSystolicPE_257_io_clear_o_d;
  wire                uSystolicPE_257_io_ifm_sign_d;
  wire                uSystolicPE_257_io_ifm_dff_d;
  wire                uSystolicPE_257_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_257_io_randW_d;
  wire       [14:0]   uSystolicPE_257_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_257_io_ofm_d;
  wire                uSystolicPE_258_io_mac_done_d;
  wire                uSystolicPE_258_io_enable_i_d;
  wire                uSystolicPE_258_io_clear_i_d;
  wire                uSystolicPE_258_io_enable_w_d;
  wire                uSystolicPE_258_io_clear_w_d;
  wire                uSystolicPE_258_io_enable_o_d;
  wire                uSystolicPE_258_io_clear_o_d;
  wire                uSystolicPE_258_io_ifm_sign_d;
  wire                uSystolicPE_258_io_ifm_dff_d;
  wire                uSystolicPE_258_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_258_io_randW_d;
  wire       [14:0]   uSystolicPE_258_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_258_io_ofm_d;
  wire                uSystolicPE_259_io_mac_done_d;
  wire                uSystolicPE_259_io_enable_i_d;
  wire                uSystolicPE_259_io_clear_i_d;
  wire                uSystolicPE_259_io_enable_w_d;
  wire                uSystolicPE_259_io_clear_w_d;
  wire                uSystolicPE_259_io_enable_o_d;
  wire                uSystolicPE_259_io_clear_o_d;
  wire                uSystolicPE_259_io_ifm_sign_d;
  wire                uSystolicPE_259_io_ifm_dff_d;
  wire                uSystolicPE_259_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_259_io_randW_d;
  wire       [14:0]   uSystolicPE_259_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_259_io_ofm_d;
  wire                uSystolicPE_260_io_mac_done_d;
  wire                uSystolicPE_260_io_enable_i_d;
  wire                uSystolicPE_260_io_clear_i_d;
  wire                uSystolicPE_260_io_enable_w_d;
  wire                uSystolicPE_260_io_clear_w_d;
  wire                uSystolicPE_260_io_enable_o_d;
  wire                uSystolicPE_260_io_clear_o_d;
  wire                uSystolicPE_260_io_ifm_sign_d;
  wire                uSystolicPE_260_io_ifm_dff_d;
  wire                uSystolicPE_260_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_260_io_randW_d;
  wire       [14:0]   uSystolicPE_260_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_260_io_ofm_d;
  wire                uSystolicPE_261_io_mac_done_d;
  wire                uSystolicPE_261_io_enable_i_d;
  wire                uSystolicPE_261_io_clear_i_d;
  wire                uSystolicPE_261_io_enable_w_d;
  wire                uSystolicPE_261_io_clear_w_d;
  wire                uSystolicPE_261_io_enable_o_d;
  wire                uSystolicPE_261_io_clear_o_d;
  wire                uSystolicPE_261_io_ifm_sign_d;
  wire                uSystolicPE_261_io_ifm_dff_d;
  wire                uSystolicPE_261_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_261_io_randW_d;
  wire       [14:0]   uSystolicPE_261_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_261_io_ofm_d;
  wire                uSystolicPE_262_io_mac_done_d;
  wire                uSystolicPE_262_io_enable_i_d;
  wire                uSystolicPE_262_io_clear_i_d;
  wire                uSystolicPE_262_io_enable_w_d;
  wire                uSystolicPE_262_io_clear_w_d;
  wire                uSystolicPE_262_io_enable_o_d;
  wire                uSystolicPE_262_io_clear_o_d;
  wire                uSystolicPE_262_io_ifm_sign_d;
  wire                uSystolicPE_262_io_ifm_dff_d;
  wire                uSystolicPE_262_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_262_io_randW_d;
  wire       [14:0]   uSystolicPE_262_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_262_io_ofm_d;
  wire                uSystolicPE_263_io_mac_done_d;
  wire                uSystolicPE_263_io_enable_i_d;
  wire                uSystolicPE_263_io_clear_i_d;
  wire                uSystolicPE_263_io_enable_w_d;
  wire                uSystolicPE_263_io_clear_w_d;
  wire                uSystolicPE_263_io_enable_o_d;
  wire                uSystolicPE_263_io_clear_o_d;
  wire                uSystolicPE_263_io_ifm_sign_d;
  wire                uSystolicPE_263_io_ifm_dff_d;
  wire                uSystolicPE_263_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_263_io_randW_d;
  wire       [14:0]   uSystolicPE_263_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_263_io_ofm_d;
  wire                uSystolicPE_264_io_mac_done_d;
  wire                uSystolicPE_264_io_enable_i_d;
  wire                uSystolicPE_264_io_clear_i_d;
  wire                uSystolicPE_264_io_enable_w_d;
  wire                uSystolicPE_264_io_clear_w_d;
  wire                uSystolicPE_264_io_enable_o_d;
  wire                uSystolicPE_264_io_clear_o_d;
  wire                uSystolicPE_264_io_ifm_sign_d;
  wire                uSystolicPE_264_io_ifm_dff_d;
  wire                uSystolicPE_264_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_264_io_randW_d;
  wire       [14:0]   uSystolicPE_264_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_264_io_ofm_d;
  wire                uSystolicPE_265_io_mac_done_d;
  wire                uSystolicPE_265_io_enable_i_d;
  wire                uSystolicPE_265_io_clear_i_d;
  wire                uSystolicPE_265_io_enable_w_d;
  wire                uSystolicPE_265_io_clear_w_d;
  wire                uSystolicPE_265_io_enable_o_d;
  wire                uSystolicPE_265_io_clear_o_d;
  wire                uSystolicPE_265_io_ifm_sign_d;
  wire                uSystolicPE_265_io_ifm_dff_d;
  wire                uSystolicPE_265_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_265_io_randW_d;
  wire       [14:0]   uSystolicPE_265_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_265_io_ofm_d;
  wire                uSystolicPE_266_io_mac_done_d;
  wire                uSystolicPE_266_io_enable_i_d;
  wire                uSystolicPE_266_io_clear_i_d;
  wire                uSystolicPE_266_io_enable_w_d;
  wire                uSystolicPE_266_io_clear_w_d;
  wire                uSystolicPE_266_io_enable_o_d;
  wire                uSystolicPE_266_io_clear_o_d;
  wire                uSystolicPE_266_io_ifm_sign_d;
  wire                uSystolicPE_266_io_ifm_dff_d;
  wire                uSystolicPE_266_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_266_io_randW_d;
  wire       [14:0]   uSystolicPE_266_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_266_io_ofm_d;
  wire                uSystolicPE_267_io_mac_done_d;
  wire                uSystolicPE_267_io_enable_i_d;
  wire                uSystolicPE_267_io_clear_i_d;
  wire                uSystolicPE_267_io_enable_w_d;
  wire                uSystolicPE_267_io_clear_w_d;
  wire                uSystolicPE_267_io_enable_o_d;
  wire                uSystolicPE_267_io_clear_o_d;
  wire                uSystolicPE_267_io_ifm_sign_d;
  wire                uSystolicPE_267_io_ifm_dff_d;
  wire                uSystolicPE_267_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_267_io_randW_d;
  wire       [14:0]   uSystolicPE_267_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_267_io_ofm_d;
  wire                uSystolicPE_268_io_mac_done_d;
  wire                uSystolicPE_268_io_enable_i_d;
  wire                uSystolicPE_268_io_clear_i_d;
  wire                uSystolicPE_268_io_enable_w_d;
  wire                uSystolicPE_268_io_clear_w_d;
  wire                uSystolicPE_268_io_enable_o_d;
  wire                uSystolicPE_268_io_clear_o_d;
  wire                uSystolicPE_268_io_ifm_sign_d;
  wire                uSystolicPE_268_io_ifm_dff_d;
  wire                uSystolicPE_268_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_268_io_randW_d;
  wire       [14:0]   uSystolicPE_268_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_268_io_ofm_d;
  wire                uSystolicPE_269_io_mac_done_d;
  wire                uSystolicPE_269_io_enable_i_d;
  wire                uSystolicPE_269_io_clear_i_d;
  wire                uSystolicPE_269_io_enable_w_d;
  wire                uSystolicPE_269_io_clear_w_d;
  wire                uSystolicPE_269_io_enable_o_d;
  wire                uSystolicPE_269_io_clear_o_d;
  wire                uSystolicPE_269_io_ifm_sign_d;
  wire                uSystolicPE_269_io_ifm_dff_d;
  wire                uSystolicPE_269_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_269_io_randW_d;
  wire       [14:0]   uSystolicPE_269_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_269_io_ofm_d;
  wire                uSystolicPEBorder_18_io_mac_done_d;
  wire                uSystolicPEBorder_18_io_enable_i_d;
  wire                uSystolicPEBorder_18_io_clear_i_d;
  wire                uSystolicPEBorder_18_io_enable_w_d;
  wire                uSystolicPEBorder_18_io_clear_w_d;
  wire                uSystolicPEBorder_18_io_enable_o_d;
  wire                uSystolicPEBorder_18_io_clear_o_d;
  wire                uSystolicPEBorder_18_io_ifm_sign_d;
  wire                uSystolicPEBorder_18_io_ifm_dff_d;
  wire                uSystolicPEBorder_18_io_wght_sign_d;
  wire       [14:0]   uSystolicPEBorder_18_io_randW_d;
  wire       [14:0]   uSystolicPEBorder_18_io_wght_abs_d;
  wire       [31:0]   uSystolicPEBorder_18_io_ofm_d;
  wire                uSystolicPE_270_io_mac_done_d;
  wire                uSystolicPE_270_io_enable_i_d;
  wire                uSystolicPE_270_io_clear_i_d;
  wire                uSystolicPE_270_io_enable_w_d;
  wire                uSystolicPE_270_io_clear_w_d;
  wire                uSystolicPE_270_io_enable_o_d;
  wire                uSystolicPE_270_io_clear_o_d;
  wire                uSystolicPE_270_io_ifm_sign_d;
  wire                uSystolicPE_270_io_ifm_dff_d;
  wire                uSystolicPE_270_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_270_io_randW_d;
  wire       [14:0]   uSystolicPE_270_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_270_io_ofm_d;
  wire                uSystolicPE_271_io_mac_done_d;
  wire                uSystolicPE_271_io_enable_i_d;
  wire                uSystolicPE_271_io_clear_i_d;
  wire                uSystolicPE_271_io_enable_w_d;
  wire                uSystolicPE_271_io_clear_w_d;
  wire                uSystolicPE_271_io_enable_o_d;
  wire                uSystolicPE_271_io_clear_o_d;
  wire                uSystolicPE_271_io_ifm_sign_d;
  wire                uSystolicPE_271_io_ifm_dff_d;
  wire                uSystolicPE_271_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_271_io_randW_d;
  wire       [14:0]   uSystolicPE_271_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_271_io_ofm_d;
  wire                uSystolicPE_272_io_mac_done_d;
  wire                uSystolicPE_272_io_enable_i_d;
  wire                uSystolicPE_272_io_clear_i_d;
  wire                uSystolicPE_272_io_enable_w_d;
  wire                uSystolicPE_272_io_clear_w_d;
  wire                uSystolicPE_272_io_enable_o_d;
  wire                uSystolicPE_272_io_clear_o_d;
  wire                uSystolicPE_272_io_ifm_sign_d;
  wire                uSystolicPE_272_io_ifm_dff_d;
  wire                uSystolicPE_272_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_272_io_randW_d;
  wire       [14:0]   uSystolicPE_272_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_272_io_ofm_d;
  wire                uSystolicPE_273_io_mac_done_d;
  wire                uSystolicPE_273_io_enable_i_d;
  wire                uSystolicPE_273_io_clear_i_d;
  wire                uSystolicPE_273_io_enable_w_d;
  wire                uSystolicPE_273_io_clear_w_d;
  wire                uSystolicPE_273_io_enable_o_d;
  wire                uSystolicPE_273_io_clear_o_d;
  wire                uSystolicPE_273_io_ifm_sign_d;
  wire                uSystolicPE_273_io_ifm_dff_d;
  wire                uSystolicPE_273_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_273_io_randW_d;
  wire       [14:0]   uSystolicPE_273_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_273_io_ofm_d;
  wire                uSystolicPE_274_io_mac_done_d;
  wire                uSystolicPE_274_io_enable_i_d;
  wire                uSystolicPE_274_io_clear_i_d;
  wire                uSystolicPE_274_io_enable_w_d;
  wire                uSystolicPE_274_io_clear_w_d;
  wire                uSystolicPE_274_io_enable_o_d;
  wire                uSystolicPE_274_io_clear_o_d;
  wire                uSystolicPE_274_io_ifm_sign_d;
  wire                uSystolicPE_274_io_ifm_dff_d;
  wire                uSystolicPE_274_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_274_io_randW_d;
  wire       [14:0]   uSystolicPE_274_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_274_io_ofm_d;
  wire                uSystolicPE_275_io_mac_done_d;
  wire                uSystolicPE_275_io_enable_i_d;
  wire                uSystolicPE_275_io_clear_i_d;
  wire                uSystolicPE_275_io_enable_w_d;
  wire                uSystolicPE_275_io_clear_w_d;
  wire                uSystolicPE_275_io_enable_o_d;
  wire                uSystolicPE_275_io_clear_o_d;
  wire                uSystolicPE_275_io_ifm_sign_d;
  wire                uSystolicPE_275_io_ifm_dff_d;
  wire                uSystolicPE_275_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_275_io_randW_d;
  wire       [14:0]   uSystolicPE_275_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_275_io_ofm_d;
  wire                uSystolicPE_276_io_mac_done_d;
  wire                uSystolicPE_276_io_enable_i_d;
  wire                uSystolicPE_276_io_clear_i_d;
  wire                uSystolicPE_276_io_enable_w_d;
  wire                uSystolicPE_276_io_clear_w_d;
  wire                uSystolicPE_276_io_enable_o_d;
  wire                uSystolicPE_276_io_clear_o_d;
  wire                uSystolicPE_276_io_ifm_sign_d;
  wire                uSystolicPE_276_io_ifm_dff_d;
  wire                uSystolicPE_276_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_276_io_randW_d;
  wire       [14:0]   uSystolicPE_276_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_276_io_ofm_d;
  wire                uSystolicPE_277_io_mac_done_d;
  wire                uSystolicPE_277_io_enable_i_d;
  wire                uSystolicPE_277_io_clear_i_d;
  wire                uSystolicPE_277_io_enable_w_d;
  wire                uSystolicPE_277_io_clear_w_d;
  wire                uSystolicPE_277_io_enable_o_d;
  wire                uSystolicPE_277_io_clear_o_d;
  wire                uSystolicPE_277_io_ifm_sign_d;
  wire                uSystolicPE_277_io_ifm_dff_d;
  wire                uSystolicPE_277_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_277_io_randW_d;
  wire       [14:0]   uSystolicPE_277_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_277_io_ofm_d;
  wire                uSystolicPE_278_io_mac_done_d;
  wire                uSystolicPE_278_io_enable_i_d;
  wire                uSystolicPE_278_io_clear_i_d;
  wire                uSystolicPE_278_io_enable_w_d;
  wire                uSystolicPE_278_io_clear_w_d;
  wire                uSystolicPE_278_io_enable_o_d;
  wire                uSystolicPE_278_io_clear_o_d;
  wire                uSystolicPE_278_io_ifm_sign_d;
  wire                uSystolicPE_278_io_ifm_dff_d;
  wire                uSystolicPE_278_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_278_io_randW_d;
  wire       [14:0]   uSystolicPE_278_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_278_io_ofm_d;
  wire                uSystolicPE_279_io_mac_done_d;
  wire                uSystolicPE_279_io_enable_i_d;
  wire                uSystolicPE_279_io_clear_i_d;
  wire                uSystolicPE_279_io_enable_w_d;
  wire                uSystolicPE_279_io_clear_w_d;
  wire                uSystolicPE_279_io_enable_o_d;
  wire                uSystolicPE_279_io_clear_o_d;
  wire                uSystolicPE_279_io_ifm_sign_d;
  wire                uSystolicPE_279_io_ifm_dff_d;
  wire                uSystolicPE_279_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_279_io_randW_d;
  wire       [14:0]   uSystolicPE_279_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_279_io_ofm_d;
  wire                uSystolicPE_280_io_mac_done_d;
  wire                uSystolicPE_280_io_enable_i_d;
  wire                uSystolicPE_280_io_clear_i_d;
  wire                uSystolicPE_280_io_enable_w_d;
  wire                uSystolicPE_280_io_clear_w_d;
  wire                uSystolicPE_280_io_enable_o_d;
  wire                uSystolicPE_280_io_clear_o_d;
  wire                uSystolicPE_280_io_ifm_sign_d;
  wire                uSystolicPE_280_io_ifm_dff_d;
  wire                uSystolicPE_280_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_280_io_randW_d;
  wire       [14:0]   uSystolicPE_280_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_280_io_ofm_d;
  wire                uSystolicPE_281_io_mac_done_d;
  wire                uSystolicPE_281_io_enable_i_d;
  wire                uSystolicPE_281_io_clear_i_d;
  wire                uSystolicPE_281_io_enable_w_d;
  wire                uSystolicPE_281_io_clear_w_d;
  wire                uSystolicPE_281_io_enable_o_d;
  wire                uSystolicPE_281_io_clear_o_d;
  wire                uSystolicPE_281_io_ifm_sign_d;
  wire                uSystolicPE_281_io_ifm_dff_d;
  wire                uSystolicPE_281_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_281_io_randW_d;
  wire       [14:0]   uSystolicPE_281_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_281_io_ofm_d;
  wire                uSystolicPE_282_io_mac_done_d;
  wire                uSystolicPE_282_io_enable_i_d;
  wire                uSystolicPE_282_io_clear_i_d;
  wire                uSystolicPE_282_io_enable_w_d;
  wire                uSystolicPE_282_io_clear_w_d;
  wire                uSystolicPE_282_io_enable_o_d;
  wire                uSystolicPE_282_io_clear_o_d;
  wire                uSystolicPE_282_io_ifm_sign_d;
  wire                uSystolicPE_282_io_ifm_dff_d;
  wire                uSystolicPE_282_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_282_io_randW_d;
  wire       [14:0]   uSystolicPE_282_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_282_io_ofm_d;
  wire                uSystolicPE_283_io_mac_done_d;
  wire                uSystolicPE_283_io_enable_i_d;
  wire                uSystolicPE_283_io_clear_i_d;
  wire                uSystolicPE_283_io_enable_w_d;
  wire                uSystolicPE_283_io_clear_w_d;
  wire                uSystolicPE_283_io_enable_o_d;
  wire                uSystolicPE_283_io_clear_o_d;
  wire                uSystolicPE_283_io_ifm_sign_d;
  wire                uSystolicPE_283_io_ifm_dff_d;
  wire                uSystolicPE_283_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_283_io_randW_d;
  wire       [14:0]   uSystolicPE_283_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_283_io_ofm_d;
  wire                uSystolicPE_284_io_mac_done_d;
  wire                uSystolicPE_284_io_enable_i_d;
  wire                uSystolicPE_284_io_clear_i_d;
  wire                uSystolicPE_284_io_enable_w_d;
  wire                uSystolicPE_284_io_clear_w_d;
  wire                uSystolicPE_284_io_enable_o_d;
  wire                uSystolicPE_284_io_clear_o_d;
  wire                uSystolicPE_284_io_ifm_sign_d;
  wire                uSystolicPE_284_io_ifm_dff_d;
  wire                uSystolicPE_284_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_284_io_randW_d;
  wire       [14:0]   uSystolicPE_284_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_284_io_ofm_d;
  wire                uSystolicPEBorder_19_io_mac_done_d;
  wire                uSystolicPEBorder_19_io_enable_i_d;
  wire                uSystolicPEBorder_19_io_clear_i_d;
  wire                uSystolicPEBorder_19_io_enable_w_d;
  wire                uSystolicPEBorder_19_io_clear_w_d;
  wire                uSystolicPEBorder_19_io_enable_o_d;
  wire                uSystolicPEBorder_19_io_clear_o_d;
  wire                uSystolicPEBorder_19_io_ifm_sign_d;
  wire                uSystolicPEBorder_19_io_ifm_dff_d;
  wire                uSystolicPEBorder_19_io_wght_sign_d;
  wire       [14:0]   uSystolicPEBorder_19_io_randW_d;
  wire       [14:0]   uSystolicPEBorder_19_io_wght_abs_d;
  wire       [31:0]   uSystolicPEBorder_19_io_ofm_d;
  wire                uSystolicPE_285_io_mac_done_d;
  wire                uSystolicPE_285_io_enable_i_d;
  wire                uSystolicPE_285_io_clear_i_d;
  wire                uSystolicPE_285_io_enable_w_d;
  wire                uSystolicPE_285_io_clear_w_d;
  wire                uSystolicPE_285_io_enable_o_d;
  wire                uSystolicPE_285_io_clear_o_d;
  wire                uSystolicPE_285_io_ifm_sign_d;
  wire                uSystolicPE_285_io_ifm_dff_d;
  wire                uSystolicPE_285_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_285_io_randW_d;
  wire       [14:0]   uSystolicPE_285_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_285_io_ofm_d;
  wire                uSystolicPE_286_io_mac_done_d;
  wire                uSystolicPE_286_io_enable_i_d;
  wire                uSystolicPE_286_io_clear_i_d;
  wire                uSystolicPE_286_io_enable_w_d;
  wire                uSystolicPE_286_io_clear_w_d;
  wire                uSystolicPE_286_io_enable_o_d;
  wire                uSystolicPE_286_io_clear_o_d;
  wire                uSystolicPE_286_io_ifm_sign_d;
  wire                uSystolicPE_286_io_ifm_dff_d;
  wire                uSystolicPE_286_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_286_io_randW_d;
  wire       [14:0]   uSystolicPE_286_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_286_io_ofm_d;
  wire                uSystolicPE_287_io_mac_done_d;
  wire                uSystolicPE_287_io_enable_i_d;
  wire                uSystolicPE_287_io_clear_i_d;
  wire                uSystolicPE_287_io_enable_w_d;
  wire                uSystolicPE_287_io_clear_w_d;
  wire                uSystolicPE_287_io_enable_o_d;
  wire                uSystolicPE_287_io_clear_o_d;
  wire                uSystolicPE_287_io_ifm_sign_d;
  wire                uSystolicPE_287_io_ifm_dff_d;
  wire                uSystolicPE_287_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_287_io_randW_d;
  wire       [14:0]   uSystolicPE_287_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_287_io_ofm_d;
  wire                uSystolicPE_288_io_mac_done_d;
  wire                uSystolicPE_288_io_enable_i_d;
  wire                uSystolicPE_288_io_clear_i_d;
  wire                uSystolicPE_288_io_enable_w_d;
  wire                uSystolicPE_288_io_clear_w_d;
  wire                uSystolicPE_288_io_enable_o_d;
  wire                uSystolicPE_288_io_clear_o_d;
  wire                uSystolicPE_288_io_ifm_sign_d;
  wire                uSystolicPE_288_io_ifm_dff_d;
  wire                uSystolicPE_288_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_288_io_randW_d;
  wire       [14:0]   uSystolicPE_288_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_288_io_ofm_d;
  wire                uSystolicPE_289_io_mac_done_d;
  wire                uSystolicPE_289_io_enable_i_d;
  wire                uSystolicPE_289_io_clear_i_d;
  wire                uSystolicPE_289_io_enable_w_d;
  wire                uSystolicPE_289_io_clear_w_d;
  wire                uSystolicPE_289_io_enable_o_d;
  wire                uSystolicPE_289_io_clear_o_d;
  wire                uSystolicPE_289_io_ifm_sign_d;
  wire                uSystolicPE_289_io_ifm_dff_d;
  wire                uSystolicPE_289_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_289_io_randW_d;
  wire       [14:0]   uSystolicPE_289_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_289_io_ofm_d;
  wire                uSystolicPE_290_io_mac_done_d;
  wire                uSystolicPE_290_io_enable_i_d;
  wire                uSystolicPE_290_io_clear_i_d;
  wire                uSystolicPE_290_io_enable_w_d;
  wire                uSystolicPE_290_io_clear_w_d;
  wire                uSystolicPE_290_io_enable_o_d;
  wire                uSystolicPE_290_io_clear_o_d;
  wire                uSystolicPE_290_io_ifm_sign_d;
  wire                uSystolicPE_290_io_ifm_dff_d;
  wire                uSystolicPE_290_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_290_io_randW_d;
  wire       [14:0]   uSystolicPE_290_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_290_io_ofm_d;
  wire                uSystolicPE_291_io_mac_done_d;
  wire                uSystolicPE_291_io_enable_i_d;
  wire                uSystolicPE_291_io_clear_i_d;
  wire                uSystolicPE_291_io_enable_w_d;
  wire                uSystolicPE_291_io_clear_w_d;
  wire                uSystolicPE_291_io_enable_o_d;
  wire                uSystolicPE_291_io_clear_o_d;
  wire                uSystolicPE_291_io_ifm_sign_d;
  wire                uSystolicPE_291_io_ifm_dff_d;
  wire                uSystolicPE_291_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_291_io_randW_d;
  wire       [14:0]   uSystolicPE_291_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_291_io_ofm_d;
  wire                uSystolicPE_292_io_mac_done_d;
  wire                uSystolicPE_292_io_enable_i_d;
  wire                uSystolicPE_292_io_clear_i_d;
  wire                uSystolicPE_292_io_enable_w_d;
  wire                uSystolicPE_292_io_clear_w_d;
  wire                uSystolicPE_292_io_enable_o_d;
  wire                uSystolicPE_292_io_clear_o_d;
  wire                uSystolicPE_292_io_ifm_sign_d;
  wire                uSystolicPE_292_io_ifm_dff_d;
  wire                uSystolicPE_292_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_292_io_randW_d;
  wire       [14:0]   uSystolicPE_292_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_292_io_ofm_d;
  wire                uSystolicPE_293_io_mac_done_d;
  wire                uSystolicPE_293_io_enable_i_d;
  wire                uSystolicPE_293_io_clear_i_d;
  wire                uSystolicPE_293_io_enable_w_d;
  wire                uSystolicPE_293_io_clear_w_d;
  wire                uSystolicPE_293_io_enable_o_d;
  wire                uSystolicPE_293_io_clear_o_d;
  wire                uSystolicPE_293_io_ifm_sign_d;
  wire                uSystolicPE_293_io_ifm_dff_d;
  wire                uSystolicPE_293_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_293_io_randW_d;
  wire       [14:0]   uSystolicPE_293_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_293_io_ofm_d;
  wire                uSystolicPE_294_io_mac_done_d;
  wire                uSystolicPE_294_io_enable_i_d;
  wire                uSystolicPE_294_io_clear_i_d;
  wire                uSystolicPE_294_io_enable_w_d;
  wire                uSystolicPE_294_io_clear_w_d;
  wire                uSystolicPE_294_io_enable_o_d;
  wire                uSystolicPE_294_io_clear_o_d;
  wire                uSystolicPE_294_io_ifm_sign_d;
  wire                uSystolicPE_294_io_ifm_dff_d;
  wire                uSystolicPE_294_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_294_io_randW_d;
  wire       [14:0]   uSystolicPE_294_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_294_io_ofm_d;
  wire                uSystolicPE_295_io_mac_done_d;
  wire                uSystolicPE_295_io_enable_i_d;
  wire                uSystolicPE_295_io_clear_i_d;
  wire                uSystolicPE_295_io_enable_w_d;
  wire                uSystolicPE_295_io_clear_w_d;
  wire                uSystolicPE_295_io_enable_o_d;
  wire                uSystolicPE_295_io_clear_o_d;
  wire                uSystolicPE_295_io_ifm_sign_d;
  wire                uSystolicPE_295_io_ifm_dff_d;
  wire                uSystolicPE_295_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_295_io_randW_d;
  wire       [14:0]   uSystolicPE_295_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_295_io_ofm_d;
  wire                uSystolicPE_296_io_mac_done_d;
  wire                uSystolicPE_296_io_enable_i_d;
  wire                uSystolicPE_296_io_clear_i_d;
  wire                uSystolicPE_296_io_enable_w_d;
  wire                uSystolicPE_296_io_clear_w_d;
  wire                uSystolicPE_296_io_enable_o_d;
  wire                uSystolicPE_296_io_clear_o_d;
  wire                uSystolicPE_296_io_ifm_sign_d;
  wire                uSystolicPE_296_io_ifm_dff_d;
  wire                uSystolicPE_296_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_296_io_randW_d;
  wire       [14:0]   uSystolicPE_296_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_296_io_ofm_d;
  wire                uSystolicPE_297_io_mac_done_d;
  wire                uSystolicPE_297_io_enable_i_d;
  wire                uSystolicPE_297_io_clear_i_d;
  wire                uSystolicPE_297_io_enable_w_d;
  wire                uSystolicPE_297_io_clear_w_d;
  wire                uSystolicPE_297_io_enable_o_d;
  wire                uSystolicPE_297_io_clear_o_d;
  wire                uSystolicPE_297_io_ifm_sign_d;
  wire                uSystolicPE_297_io_ifm_dff_d;
  wire                uSystolicPE_297_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_297_io_randW_d;
  wire       [14:0]   uSystolicPE_297_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_297_io_ofm_d;
  wire                uSystolicPE_298_io_mac_done_d;
  wire                uSystolicPE_298_io_enable_i_d;
  wire                uSystolicPE_298_io_clear_i_d;
  wire                uSystolicPE_298_io_enable_w_d;
  wire                uSystolicPE_298_io_clear_w_d;
  wire                uSystolicPE_298_io_enable_o_d;
  wire                uSystolicPE_298_io_clear_o_d;
  wire                uSystolicPE_298_io_ifm_sign_d;
  wire                uSystolicPE_298_io_ifm_dff_d;
  wire                uSystolicPE_298_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_298_io_randW_d;
  wire       [14:0]   uSystolicPE_298_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_298_io_ofm_d;
  wire                uSystolicPE_299_io_mac_done_d;
  wire                uSystolicPE_299_io_enable_i_d;
  wire                uSystolicPE_299_io_clear_i_d;
  wire                uSystolicPE_299_io_enable_w_d;
  wire                uSystolicPE_299_io_clear_w_d;
  wire                uSystolicPE_299_io_enable_o_d;
  wire                uSystolicPE_299_io_clear_o_d;
  wire                uSystolicPE_299_io_ifm_sign_d;
  wire                uSystolicPE_299_io_ifm_dff_d;
  wire                uSystolicPE_299_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_299_io_randW_d;
  wire       [14:0]   uSystolicPE_299_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_299_io_ofm_d;
  wire                uSystolicPEBorder_20_io_mac_done_d;
  wire                uSystolicPEBorder_20_io_enable_i_d;
  wire                uSystolicPEBorder_20_io_clear_i_d;
  wire                uSystolicPEBorder_20_io_enable_w_d;
  wire                uSystolicPEBorder_20_io_clear_w_d;
  wire                uSystolicPEBorder_20_io_enable_o_d;
  wire                uSystolicPEBorder_20_io_clear_o_d;
  wire                uSystolicPEBorder_20_io_ifm_sign_d;
  wire                uSystolicPEBorder_20_io_ifm_dff_d;
  wire                uSystolicPEBorder_20_io_wght_sign_d;
  wire       [14:0]   uSystolicPEBorder_20_io_randW_d;
  wire       [14:0]   uSystolicPEBorder_20_io_wght_abs_d;
  wire       [31:0]   uSystolicPEBorder_20_io_ofm_d;
  wire                uSystolicPE_300_io_mac_done_d;
  wire                uSystolicPE_300_io_enable_i_d;
  wire                uSystolicPE_300_io_clear_i_d;
  wire                uSystolicPE_300_io_enable_w_d;
  wire                uSystolicPE_300_io_clear_w_d;
  wire                uSystolicPE_300_io_enable_o_d;
  wire                uSystolicPE_300_io_clear_o_d;
  wire                uSystolicPE_300_io_ifm_sign_d;
  wire                uSystolicPE_300_io_ifm_dff_d;
  wire                uSystolicPE_300_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_300_io_randW_d;
  wire       [14:0]   uSystolicPE_300_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_300_io_ofm_d;
  wire                uSystolicPE_301_io_mac_done_d;
  wire                uSystolicPE_301_io_enable_i_d;
  wire                uSystolicPE_301_io_clear_i_d;
  wire                uSystolicPE_301_io_enable_w_d;
  wire                uSystolicPE_301_io_clear_w_d;
  wire                uSystolicPE_301_io_enable_o_d;
  wire                uSystolicPE_301_io_clear_o_d;
  wire                uSystolicPE_301_io_ifm_sign_d;
  wire                uSystolicPE_301_io_ifm_dff_d;
  wire                uSystolicPE_301_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_301_io_randW_d;
  wire       [14:0]   uSystolicPE_301_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_301_io_ofm_d;
  wire                uSystolicPE_302_io_mac_done_d;
  wire                uSystolicPE_302_io_enable_i_d;
  wire                uSystolicPE_302_io_clear_i_d;
  wire                uSystolicPE_302_io_enable_w_d;
  wire                uSystolicPE_302_io_clear_w_d;
  wire                uSystolicPE_302_io_enable_o_d;
  wire                uSystolicPE_302_io_clear_o_d;
  wire                uSystolicPE_302_io_ifm_sign_d;
  wire                uSystolicPE_302_io_ifm_dff_d;
  wire                uSystolicPE_302_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_302_io_randW_d;
  wire       [14:0]   uSystolicPE_302_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_302_io_ofm_d;
  wire                uSystolicPE_303_io_mac_done_d;
  wire                uSystolicPE_303_io_enable_i_d;
  wire                uSystolicPE_303_io_clear_i_d;
  wire                uSystolicPE_303_io_enable_w_d;
  wire                uSystolicPE_303_io_clear_w_d;
  wire                uSystolicPE_303_io_enable_o_d;
  wire                uSystolicPE_303_io_clear_o_d;
  wire                uSystolicPE_303_io_ifm_sign_d;
  wire                uSystolicPE_303_io_ifm_dff_d;
  wire                uSystolicPE_303_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_303_io_randW_d;
  wire       [14:0]   uSystolicPE_303_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_303_io_ofm_d;
  wire                uSystolicPE_304_io_mac_done_d;
  wire                uSystolicPE_304_io_enable_i_d;
  wire                uSystolicPE_304_io_clear_i_d;
  wire                uSystolicPE_304_io_enable_w_d;
  wire                uSystolicPE_304_io_clear_w_d;
  wire                uSystolicPE_304_io_enable_o_d;
  wire                uSystolicPE_304_io_clear_o_d;
  wire                uSystolicPE_304_io_ifm_sign_d;
  wire                uSystolicPE_304_io_ifm_dff_d;
  wire                uSystolicPE_304_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_304_io_randW_d;
  wire       [14:0]   uSystolicPE_304_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_304_io_ofm_d;
  wire                uSystolicPE_305_io_mac_done_d;
  wire                uSystolicPE_305_io_enable_i_d;
  wire                uSystolicPE_305_io_clear_i_d;
  wire                uSystolicPE_305_io_enable_w_d;
  wire                uSystolicPE_305_io_clear_w_d;
  wire                uSystolicPE_305_io_enable_o_d;
  wire                uSystolicPE_305_io_clear_o_d;
  wire                uSystolicPE_305_io_ifm_sign_d;
  wire                uSystolicPE_305_io_ifm_dff_d;
  wire                uSystolicPE_305_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_305_io_randW_d;
  wire       [14:0]   uSystolicPE_305_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_305_io_ofm_d;
  wire                uSystolicPE_306_io_mac_done_d;
  wire                uSystolicPE_306_io_enable_i_d;
  wire                uSystolicPE_306_io_clear_i_d;
  wire                uSystolicPE_306_io_enable_w_d;
  wire                uSystolicPE_306_io_clear_w_d;
  wire                uSystolicPE_306_io_enable_o_d;
  wire                uSystolicPE_306_io_clear_o_d;
  wire                uSystolicPE_306_io_ifm_sign_d;
  wire                uSystolicPE_306_io_ifm_dff_d;
  wire                uSystolicPE_306_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_306_io_randW_d;
  wire       [14:0]   uSystolicPE_306_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_306_io_ofm_d;
  wire                uSystolicPE_307_io_mac_done_d;
  wire                uSystolicPE_307_io_enable_i_d;
  wire                uSystolicPE_307_io_clear_i_d;
  wire                uSystolicPE_307_io_enable_w_d;
  wire                uSystolicPE_307_io_clear_w_d;
  wire                uSystolicPE_307_io_enable_o_d;
  wire                uSystolicPE_307_io_clear_o_d;
  wire                uSystolicPE_307_io_ifm_sign_d;
  wire                uSystolicPE_307_io_ifm_dff_d;
  wire                uSystolicPE_307_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_307_io_randW_d;
  wire       [14:0]   uSystolicPE_307_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_307_io_ofm_d;
  wire                uSystolicPE_308_io_mac_done_d;
  wire                uSystolicPE_308_io_enable_i_d;
  wire                uSystolicPE_308_io_clear_i_d;
  wire                uSystolicPE_308_io_enable_w_d;
  wire                uSystolicPE_308_io_clear_w_d;
  wire                uSystolicPE_308_io_enable_o_d;
  wire                uSystolicPE_308_io_clear_o_d;
  wire                uSystolicPE_308_io_ifm_sign_d;
  wire                uSystolicPE_308_io_ifm_dff_d;
  wire                uSystolicPE_308_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_308_io_randW_d;
  wire       [14:0]   uSystolicPE_308_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_308_io_ofm_d;
  wire                uSystolicPE_309_io_mac_done_d;
  wire                uSystolicPE_309_io_enable_i_d;
  wire                uSystolicPE_309_io_clear_i_d;
  wire                uSystolicPE_309_io_enable_w_d;
  wire                uSystolicPE_309_io_clear_w_d;
  wire                uSystolicPE_309_io_enable_o_d;
  wire                uSystolicPE_309_io_clear_o_d;
  wire                uSystolicPE_309_io_ifm_sign_d;
  wire                uSystolicPE_309_io_ifm_dff_d;
  wire                uSystolicPE_309_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_309_io_randW_d;
  wire       [14:0]   uSystolicPE_309_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_309_io_ofm_d;
  wire                uSystolicPE_310_io_mac_done_d;
  wire                uSystolicPE_310_io_enable_i_d;
  wire                uSystolicPE_310_io_clear_i_d;
  wire                uSystolicPE_310_io_enable_w_d;
  wire                uSystolicPE_310_io_clear_w_d;
  wire                uSystolicPE_310_io_enable_o_d;
  wire                uSystolicPE_310_io_clear_o_d;
  wire                uSystolicPE_310_io_ifm_sign_d;
  wire                uSystolicPE_310_io_ifm_dff_d;
  wire                uSystolicPE_310_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_310_io_randW_d;
  wire       [14:0]   uSystolicPE_310_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_310_io_ofm_d;
  wire                uSystolicPE_311_io_mac_done_d;
  wire                uSystolicPE_311_io_enable_i_d;
  wire                uSystolicPE_311_io_clear_i_d;
  wire                uSystolicPE_311_io_enable_w_d;
  wire                uSystolicPE_311_io_clear_w_d;
  wire                uSystolicPE_311_io_enable_o_d;
  wire                uSystolicPE_311_io_clear_o_d;
  wire                uSystolicPE_311_io_ifm_sign_d;
  wire                uSystolicPE_311_io_ifm_dff_d;
  wire                uSystolicPE_311_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_311_io_randW_d;
  wire       [14:0]   uSystolicPE_311_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_311_io_ofm_d;
  wire                uSystolicPE_312_io_mac_done_d;
  wire                uSystolicPE_312_io_enable_i_d;
  wire                uSystolicPE_312_io_clear_i_d;
  wire                uSystolicPE_312_io_enable_w_d;
  wire                uSystolicPE_312_io_clear_w_d;
  wire                uSystolicPE_312_io_enable_o_d;
  wire                uSystolicPE_312_io_clear_o_d;
  wire                uSystolicPE_312_io_ifm_sign_d;
  wire                uSystolicPE_312_io_ifm_dff_d;
  wire                uSystolicPE_312_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_312_io_randW_d;
  wire       [14:0]   uSystolicPE_312_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_312_io_ofm_d;
  wire                uSystolicPE_313_io_mac_done_d;
  wire                uSystolicPE_313_io_enable_i_d;
  wire                uSystolicPE_313_io_clear_i_d;
  wire                uSystolicPE_313_io_enable_w_d;
  wire                uSystolicPE_313_io_clear_w_d;
  wire                uSystolicPE_313_io_enable_o_d;
  wire                uSystolicPE_313_io_clear_o_d;
  wire                uSystolicPE_313_io_ifm_sign_d;
  wire                uSystolicPE_313_io_ifm_dff_d;
  wire                uSystolicPE_313_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_313_io_randW_d;
  wire       [14:0]   uSystolicPE_313_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_313_io_ofm_d;
  wire                uSystolicPE_314_io_mac_done_d;
  wire                uSystolicPE_314_io_enable_i_d;
  wire                uSystolicPE_314_io_clear_i_d;
  wire                uSystolicPE_314_io_enable_w_d;
  wire                uSystolicPE_314_io_clear_w_d;
  wire                uSystolicPE_314_io_enable_o_d;
  wire                uSystolicPE_314_io_clear_o_d;
  wire                uSystolicPE_314_io_ifm_sign_d;
  wire                uSystolicPE_314_io_ifm_dff_d;
  wire                uSystolicPE_314_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_314_io_randW_d;
  wire       [14:0]   uSystolicPE_314_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_314_io_ofm_d;
  wire                uSystolicPEBorder_21_io_mac_done_d;
  wire                uSystolicPEBorder_21_io_enable_i_d;
  wire                uSystolicPEBorder_21_io_clear_i_d;
  wire                uSystolicPEBorder_21_io_enable_w_d;
  wire                uSystolicPEBorder_21_io_clear_w_d;
  wire                uSystolicPEBorder_21_io_enable_o_d;
  wire                uSystolicPEBorder_21_io_clear_o_d;
  wire                uSystolicPEBorder_21_io_ifm_sign_d;
  wire                uSystolicPEBorder_21_io_ifm_dff_d;
  wire                uSystolicPEBorder_21_io_wght_sign_d;
  wire       [14:0]   uSystolicPEBorder_21_io_randW_d;
  wire       [14:0]   uSystolicPEBorder_21_io_wght_abs_d;
  wire       [31:0]   uSystolicPEBorder_21_io_ofm_d;
  wire                uSystolicPE_315_io_mac_done_d;
  wire                uSystolicPE_315_io_enable_i_d;
  wire                uSystolicPE_315_io_clear_i_d;
  wire                uSystolicPE_315_io_enable_w_d;
  wire                uSystolicPE_315_io_clear_w_d;
  wire                uSystolicPE_315_io_enable_o_d;
  wire                uSystolicPE_315_io_clear_o_d;
  wire                uSystolicPE_315_io_ifm_sign_d;
  wire                uSystolicPE_315_io_ifm_dff_d;
  wire                uSystolicPE_315_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_315_io_randW_d;
  wire       [14:0]   uSystolicPE_315_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_315_io_ofm_d;
  wire                uSystolicPE_316_io_mac_done_d;
  wire                uSystolicPE_316_io_enable_i_d;
  wire                uSystolicPE_316_io_clear_i_d;
  wire                uSystolicPE_316_io_enable_w_d;
  wire                uSystolicPE_316_io_clear_w_d;
  wire                uSystolicPE_316_io_enable_o_d;
  wire                uSystolicPE_316_io_clear_o_d;
  wire                uSystolicPE_316_io_ifm_sign_d;
  wire                uSystolicPE_316_io_ifm_dff_d;
  wire                uSystolicPE_316_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_316_io_randW_d;
  wire       [14:0]   uSystolicPE_316_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_316_io_ofm_d;
  wire                uSystolicPE_317_io_mac_done_d;
  wire                uSystolicPE_317_io_enable_i_d;
  wire                uSystolicPE_317_io_clear_i_d;
  wire                uSystolicPE_317_io_enable_w_d;
  wire                uSystolicPE_317_io_clear_w_d;
  wire                uSystolicPE_317_io_enable_o_d;
  wire                uSystolicPE_317_io_clear_o_d;
  wire                uSystolicPE_317_io_ifm_sign_d;
  wire                uSystolicPE_317_io_ifm_dff_d;
  wire                uSystolicPE_317_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_317_io_randW_d;
  wire       [14:0]   uSystolicPE_317_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_317_io_ofm_d;
  wire                uSystolicPE_318_io_mac_done_d;
  wire                uSystolicPE_318_io_enable_i_d;
  wire                uSystolicPE_318_io_clear_i_d;
  wire                uSystolicPE_318_io_enable_w_d;
  wire                uSystolicPE_318_io_clear_w_d;
  wire                uSystolicPE_318_io_enable_o_d;
  wire                uSystolicPE_318_io_clear_o_d;
  wire                uSystolicPE_318_io_ifm_sign_d;
  wire                uSystolicPE_318_io_ifm_dff_d;
  wire                uSystolicPE_318_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_318_io_randW_d;
  wire       [14:0]   uSystolicPE_318_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_318_io_ofm_d;
  wire                uSystolicPE_319_io_mac_done_d;
  wire                uSystolicPE_319_io_enable_i_d;
  wire                uSystolicPE_319_io_clear_i_d;
  wire                uSystolicPE_319_io_enable_w_d;
  wire                uSystolicPE_319_io_clear_w_d;
  wire                uSystolicPE_319_io_enable_o_d;
  wire                uSystolicPE_319_io_clear_o_d;
  wire                uSystolicPE_319_io_ifm_sign_d;
  wire                uSystolicPE_319_io_ifm_dff_d;
  wire                uSystolicPE_319_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_319_io_randW_d;
  wire       [14:0]   uSystolicPE_319_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_319_io_ofm_d;
  wire                uSystolicPE_320_io_mac_done_d;
  wire                uSystolicPE_320_io_enable_i_d;
  wire                uSystolicPE_320_io_clear_i_d;
  wire                uSystolicPE_320_io_enable_w_d;
  wire                uSystolicPE_320_io_clear_w_d;
  wire                uSystolicPE_320_io_enable_o_d;
  wire                uSystolicPE_320_io_clear_o_d;
  wire                uSystolicPE_320_io_ifm_sign_d;
  wire                uSystolicPE_320_io_ifm_dff_d;
  wire                uSystolicPE_320_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_320_io_randW_d;
  wire       [14:0]   uSystolicPE_320_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_320_io_ofm_d;
  wire                uSystolicPE_321_io_mac_done_d;
  wire                uSystolicPE_321_io_enable_i_d;
  wire                uSystolicPE_321_io_clear_i_d;
  wire                uSystolicPE_321_io_enable_w_d;
  wire                uSystolicPE_321_io_clear_w_d;
  wire                uSystolicPE_321_io_enable_o_d;
  wire                uSystolicPE_321_io_clear_o_d;
  wire                uSystolicPE_321_io_ifm_sign_d;
  wire                uSystolicPE_321_io_ifm_dff_d;
  wire                uSystolicPE_321_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_321_io_randW_d;
  wire       [14:0]   uSystolicPE_321_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_321_io_ofm_d;
  wire                uSystolicPE_322_io_mac_done_d;
  wire                uSystolicPE_322_io_enable_i_d;
  wire                uSystolicPE_322_io_clear_i_d;
  wire                uSystolicPE_322_io_enable_w_d;
  wire                uSystolicPE_322_io_clear_w_d;
  wire                uSystolicPE_322_io_enable_o_d;
  wire                uSystolicPE_322_io_clear_o_d;
  wire                uSystolicPE_322_io_ifm_sign_d;
  wire                uSystolicPE_322_io_ifm_dff_d;
  wire                uSystolicPE_322_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_322_io_randW_d;
  wire       [14:0]   uSystolicPE_322_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_322_io_ofm_d;
  wire                uSystolicPE_323_io_mac_done_d;
  wire                uSystolicPE_323_io_enable_i_d;
  wire                uSystolicPE_323_io_clear_i_d;
  wire                uSystolicPE_323_io_enable_w_d;
  wire                uSystolicPE_323_io_clear_w_d;
  wire                uSystolicPE_323_io_enable_o_d;
  wire                uSystolicPE_323_io_clear_o_d;
  wire                uSystolicPE_323_io_ifm_sign_d;
  wire                uSystolicPE_323_io_ifm_dff_d;
  wire                uSystolicPE_323_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_323_io_randW_d;
  wire       [14:0]   uSystolicPE_323_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_323_io_ofm_d;
  wire                uSystolicPE_324_io_mac_done_d;
  wire                uSystolicPE_324_io_enable_i_d;
  wire                uSystolicPE_324_io_clear_i_d;
  wire                uSystolicPE_324_io_enable_w_d;
  wire                uSystolicPE_324_io_clear_w_d;
  wire                uSystolicPE_324_io_enable_o_d;
  wire                uSystolicPE_324_io_clear_o_d;
  wire                uSystolicPE_324_io_ifm_sign_d;
  wire                uSystolicPE_324_io_ifm_dff_d;
  wire                uSystolicPE_324_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_324_io_randW_d;
  wire       [14:0]   uSystolicPE_324_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_324_io_ofm_d;
  wire                uSystolicPE_325_io_mac_done_d;
  wire                uSystolicPE_325_io_enable_i_d;
  wire                uSystolicPE_325_io_clear_i_d;
  wire                uSystolicPE_325_io_enable_w_d;
  wire                uSystolicPE_325_io_clear_w_d;
  wire                uSystolicPE_325_io_enable_o_d;
  wire                uSystolicPE_325_io_clear_o_d;
  wire                uSystolicPE_325_io_ifm_sign_d;
  wire                uSystolicPE_325_io_ifm_dff_d;
  wire                uSystolicPE_325_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_325_io_randW_d;
  wire       [14:0]   uSystolicPE_325_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_325_io_ofm_d;
  wire                uSystolicPE_326_io_mac_done_d;
  wire                uSystolicPE_326_io_enable_i_d;
  wire                uSystolicPE_326_io_clear_i_d;
  wire                uSystolicPE_326_io_enable_w_d;
  wire                uSystolicPE_326_io_clear_w_d;
  wire                uSystolicPE_326_io_enable_o_d;
  wire                uSystolicPE_326_io_clear_o_d;
  wire                uSystolicPE_326_io_ifm_sign_d;
  wire                uSystolicPE_326_io_ifm_dff_d;
  wire                uSystolicPE_326_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_326_io_randW_d;
  wire       [14:0]   uSystolicPE_326_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_326_io_ofm_d;
  wire                uSystolicPE_327_io_mac_done_d;
  wire                uSystolicPE_327_io_enable_i_d;
  wire                uSystolicPE_327_io_clear_i_d;
  wire                uSystolicPE_327_io_enable_w_d;
  wire                uSystolicPE_327_io_clear_w_d;
  wire                uSystolicPE_327_io_enable_o_d;
  wire                uSystolicPE_327_io_clear_o_d;
  wire                uSystolicPE_327_io_ifm_sign_d;
  wire                uSystolicPE_327_io_ifm_dff_d;
  wire                uSystolicPE_327_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_327_io_randW_d;
  wire       [14:0]   uSystolicPE_327_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_327_io_ofm_d;
  wire                uSystolicPE_328_io_mac_done_d;
  wire                uSystolicPE_328_io_enable_i_d;
  wire                uSystolicPE_328_io_clear_i_d;
  wire                uSystolicPE_328_io_enable_w_d;
  wire                uSystolicPE_328_io_clear_w_d;
  wire                uSystolicPE_328_io_enable_o_d;
  wire                uSystolicPE_328_io_clear_o_d;
  wire                uSystolicPE_328_io_ifm_sign_d;
  wire                uSystolicPE_328_io_ifm_dff_d;
  wire                uSystolicPE_328_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_328_io_randW_d;
  wire       [14:0]   uSystolicPE_328_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_328_io_ofm_d;
  wire                uSystolicPE_329_io_mac_done_d;
  wire                uSystolicPE_329_io_enable_i_d;
  wire                uSystolicPE_329_io_clear_i_d;
  wire                uSystolicPE_329_io_enable_w_d;
  wire                uSystolicPE_329_io_clear_w_d;
  wire                uSystolicPE_329_io_enable_o_d;
  wire                uSystolicPE_329_io_clear_o_d;
  wire                uSystolicPE_329_io_ifm_sign_d;
  wire                uSystolicPE_329_io_ifm_dff_d;
  wire                uSystolicPE_329_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_329_io_randW_d;
  wire       [14:0]   uSystolicPE_329_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_329_io_ofm_d;
  wire                uSystolicPEBorder_22_io_mac_done_d;
  wire                uSystolicPEBorder_22_io_enable_i_d;
  wire                uSystolicPEBorder_22_io_clear_i_d;
  wire                uSystolicPEBorder_22_io_enable_w_d;
  wire                uSystolicPEBorder_22_io_clear_w_d;
  wire                uSystolicPEBorder_22_io_enable_o_d;
  wire                uSystolicPEBorder_22_io_clear_o_d;
  wire                uSystolicPEBorder_22_io_ifm_sign_d;
  wire                uSystolicPEBorder_22_io_ifm_dff_d;
  wire                uSystolicPEBorder_22_io_wght_sign_d;
  wire       [14:0]   uSystolicPEBorder_22_io_randW_d;
  wire       [14:0]   uSystolicPEBorder_22_io_wght_abs_d;
  wire       [31:0]   uSystolicPEBorder_22_io_ofm_d;
  wire                uSystolicPE_330_io_mac_done_d;
  wire                uSystolicPE_330_io_enable_i_d;
  wire                uSystolicPE_330_io_clear_i_d;
  wire                uSystolicPE_330_io_enable_w_d;
  wire                uSystolicPE_330_io_clear_w_d;
  wire                uSystolicPE_330_io_enable_o_d;
  wire                uSystolicPE_330_io_clear_o_d;
  wire                uSystolicPE_330_io_ifm_sign_d;
  wire                uSystolicPE_330_io_ifm_dff_d;
  wire                uSystolicPE_330_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_330_io_randW_d;
  wire       [14:0]   uSystolicPE_330_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_330_io_ofm_d;
  wire                uSystolicPE_331_io_mac_done_d;
  wire                uSystolicPE_331_io_enable_i_d;
  wire                uSystolicPE_331_io_clear_i_d;
  wire                uSystolicPE_331_io_enable_w_d;
  wire                uSystolicPE_331_io_clear_w_d;
  wire                uSystolicPE_331_io_enable_o_d;
  wire                uSystolicPE_331_io_clear_o_d;
  wire                uSystolicPE_331_io_ifm_sign_d;
  wire                uSystolicPE_331_io_ifm_dff_d;
  wire                uSystolicPE_331_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_331_io_randW_d;
  wire       [14:0]   uSystolicPE_331_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_331_io_ofm_d;
  wire                uSystolicPE_332_io_mac_done_d;
  wire                uSystolicPE_332_io_enable_i_d;
  wire                uSystolicPE_332_io_clear_i_d;
  wire                uSystolicPE_332_io_enable_w_d;
  wire                uSystolicPE_332_io_clear_w_d;
  wire                uSystolicPE_332_io_enable_o_d;
  wire                uSystolicPE_332_io_clear_o_d;
  wire                uSystolicPE_332_io_ifm_sign_d;
  wire                uSystolicPE_332_io_ifm_dff_d;
  wire                uSystolicPE_332_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_332_io_randW_d;
  wire       [14:0]   uSystolicPE_332_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_332_io_ofm_d;
  wire                uSystolicPE_333_io_mac_done_d;
  wire                uSystolicPE_333_io_enable_i_d;
  wire                uSystolicPE_333_io_clear_i_d;
  wire                uSystolicPE_333_io_enable_w_d;
  wire                uSystolicPE_333_io_clear_w_d;
  wire                uSystolicPE_333_io_enable_o_d;
  wire                uSystolicPE_333_io_clear_o_d;
  wire                uSystolicPE_333_io_ifm_sign_d;
  wire                uSystolicPE_333_io_ifm_dff_d;
  wire                uSystolicPE_333_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_333_io_randW_d;
  wire       [14:0]   uSystolicPE_333_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_333_io_ofm_d;
  wire                uSystolicPE_334_io_mac_done_d;
  wire                uSystolicPE_334_io_enable_i_d;
  wire                uSystolicPE_334_io_clear_i_d;
  wire                uSystolicPE_334_io_enable_w_d;
  wire                uSystolicPE_334_io_clear_w_d;
  wire                uSystolicPE_334_io_enable_o_d;
  wire                uSystolicPE_334_io_clear_o_d;
  wire                uSystolicPE_334_io_ifm_sign_d;
  wire                uSystolicPE_334_io_ifm_dff_d;
  wire                uSystolicPE_334_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_334_io_randW_d;
  wire       [14:0]   uSystolicPE_334_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_334_io_ofm_d;
  wire                uSystolicPE_335_io_mac_done_d;
  wire                uSystolicPE_335_io_enable_i_d;
  wire                uSystolicPE_335_io_clear_i_d;
  wire                uSystolicPE_335_io_enable_w_d;
  wire                uSystolicPE_335_io_clear_w_d;
  wire                uSystolicPE_335_io_enable_o_d;
  wire                uSystolicPE_335_io_clear_o_d;
  wire                uSystolicPE_335_io_ifm_sign_d;
  wire                uSystolicPE_335_io_ifm_dff_d;
  wire                uSystolicPE_335_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_335_io_randW_d;
  wire       [14:0]   uSystolicPE_335_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_335_io_ofm_d;
  wire                uSystolicPE_336_io_mac_done_d;
  wire                uSystolicPE_336_io_enable_i_d;
  wire                uSystolicPE_336_io_clear_i_d;
  wire                uSystolicPE_336_io_enable_w_d;
  wire                uSystolicPE_336_io_clear_w_d;
  wire                uSystolicPE_336_io_enable_o_d;
  wire                uSystolicPE_336_io_clear_o_d;
  wire                uSystolicPE_336_io_ifm_sign_d;
  wire                uSystolicPE_336_io_ifm_dff_d;
  wire                uSystolicPE_336_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_336_io_randW_d;
  wire       [14:0]   uSystolicPE_336_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_336_io_ofm_d;
  wire                uSystolicPE_337_io_mac_done_d;
  wire                uSystolicPE_337_io_enable_i_d;
  wire                uSystolicPE_337_io_clear_i_d;
  wire                uSystolicPE_337_io_enable_w_d;
  wire                uSystolicPE_337_io_clear_w_d;
  wire                uSystolicPE_337_io_enable_o_d;
  wire                uSystolicPE_337_io_clear_o_d;
  wire                uSystolicPE_337_io_ifm_sign_d;
  wire                uSystolicPE_337_io_ifm_dff_d;
  wire                uSystolicPE_337_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_337_io_randW_d;
  wire       [14:0]   uSystolicPE_337_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_337_io_ofm_d;
  wire                uSystolicPE_338_io_mac_done_d;
  wire                uSystolicPE_338_io_enable_i_d;
  wire                uSystolicPE_338_io_clear_i_d;
  wire                uSystolicPE_338_io_enable_w_d;
  wire                uSystolicPE_338_io_clear_w_d;
  wire                uSystolicPE_338_io_enable_o_d;
  wire                uSystolicPE_338_io_clear_o_d;
  wire                uSystolicPE_338_io_ifm_sign_d;
  wire                uSystolicPE_338_io_ifm_dff_d;
  wire                uSystolicPE_338_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_338_io_randW_d;
  wire       [14:0]   uSystolicPE_338_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_338_io_ofm_d;
  wire                uSystolicPE_339_io_mac_done_d;
  wire                uSystolicPE_339_io_enable_i_d;
  wire                uSystolicPE_339_io_clear_i_d;
  wire                uSystolicPE_339_io_enable_w_d;
  wire                uSystolicPE_339_io_clear_w_d;
  wire                uSystolicPE_339_io_enable_o_d;
  wire                uSystolicPE_339_io_clear_o_d;
  wire                uSystolicPE_339_io_ifm_sign_d;
  wire                uSystolicPE_339_io_ifm_dff_d;
  wire                uSystolicPE_339_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_339_io_randW_d;
  wire       [14:0]   uSystolicPE_339_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_339_io_ofm_d;
  wire                uSystolicPE_340_io_mac_done_d;
  wire                uSystolicPE_340_io_enable_i_d;
  wire                uSystolicPE_340_io_clear_i_d;
  wire                uSystolicPE_340_io_enable_w_d;
  wire                uSystolicPE_340_io_clear_w_d;
  wire                uSystolicPE_340_io_enable_o_d;
  wire                uSystolicPE_340_io_clear_o_d;
  wire                uSystolicPE_340_io_ifm_sign_d;
  wire                uSystolicPE_340_io_ifm_dff_d;
  wire                uSystolicPE_340_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_340_io_randW_d;
  wire       [14:0]   uSystolicPE_340_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_340_io_ofm_d;
  wire                uSystolicPE_341_io_mac_done_d;
  wire                uSystolicPE_341_io_enable_i_d;
  wire                uSystolicPE_341_io_clear_i_d;
  wire                uSystolicPE_341_io_enable_w_d;
  wire                uSystolicPE_341_io_clear_w_d;
  wire                uSystolicPE_341_io_enable_o_d;
  wire                uSystolicPE_341_io_clear_o_d;
  wire                uSystolicPE_341_io_ifm_sign_d;
  wire                uSystolicPE_341_io_ifm_dff_d;
  wire                uSystolicPE_341_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_341_io_randW_d;
  wire       [14:0]   uSystolicPE_341_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_341_io_ofm_d;
  wire                uSystolicPE_342_io_mac_done_d;
  wire                uSystolicPE_342_io_enable_i_d;
  wire                uSystolicPE_342_io_clear_i_d;
  wire                uSystolicPE_342_io_enable_w_d;
  wire                uSystolicPE_342_io_clear_w_d;
  wire                uSystolicPE_342_io_enable_o_d;
  wire                uSystolicPE_342_io_clear_o_d;
  wire                uSystolicPE_342_io_ifm_sign_d;
  wire                uSystolicPE_342_io_ifm_dff_d;
  wire                uSystolicPE_342_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_342_io_randW_d;
  wire       [14:0]   uSystolicPE_342_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_342_io_ofm_d;
  wire                uSystolicPE_343_io_mac_done_d;
  wire                uSystolicPE_343_io_enable_i_d;
  wire                uSystolicPE_343_io_clear_i_d;
  wire                uSystolicPE_343_io_enable_w_d;
  wire                uSystolicPE_343_io_clear_w_d;
  wire                uSystolicPE_343_io_enable_o_d;
  wire                uSystolicPE_343_io_clear_o_d;
  wire                uSystolicPE_343_io_ifm_sign_d;
  wire                uSystolicPE_343_io_ifm_dff_d;
  wire                uSystolicPE_343_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_343_io_randW_d;
  wire       [14:0]   uSystolicPE_343_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_343_io_ofm_d;
  wire                uSystolicPE_344_io_mac_done_d;
  wire                uSystolicPE_344_io_enable_i_d;
  wire                uSystolicPE_344_io_clear_i_d;
  wire                uSystolicPE_344_io_enable_w_d;
  wire                uSystolicPE_344_io_clear_w_d;
  wire                uSystolicPE_344_io_enable_o_d;
  wire                uSystolicPE_344_io_clear_o_d;
  wire                uSystolicPE_344_io_ifm_sign_d;
  wire                uSystolicPE_344_io_ifm_dff_d;
  wire                uSystolicPE_344_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_344_io_randW_d;
  wire       [14:0]   uSystolicPE_344_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_344_io_ofm_d;
  wire                uSystolicPEBorder_23_io_mac_done_d;
  wire                uSystolicPEBorder_23_io_enable_i_d;
  wire                uSystolicPEBorder_23_io_clear_i_d;
  wire                uSystolicPEBorder_23_io_enable_w_d;
  wire                uSystolicPEBorder_23_io_clear_w_d;
  wire                uSystolicPEBorder_23_io_enable_o_d;
  wire                uSystolicPEBorder_23_io_clear_o_d;
  wire                uSystolicPEBorder_23_io_ifm_sign_d;
  wire                uSystolicPEBorder_23_io_ifm_dff_d;
  wire                uSystolicPEBorder_23_io_wght_sign_d;
  wire       [14:0]   uSystolicPEBorder_23_io_randW_d;
  wire       [14:0]   uSystolicPEBorder_23_io_wght_abs_d;
  wire       [31:0]   uSystolicPEBorder_23_io_ofm_d;
  wire                uSystolicPE_345_io_mac_done_d;
  wire                uSystolicPE_345_io_enable_i_d;
  wire                uSystolicPE_345_io_clear_i_d;
  wire                uSystolicPE_345_io_enable_w_d;
  wire                uSystolicPE_345_io_clear_w_d;
  wire                uSystolicPE_345_io_enable_o_d;
  wire                uSystolicPE_345_io_clear_o_d;
  wire                uSystolicPE_345_io_ifm_sign_d;
  wire                uSystolicPE_345_io_ifm_dff_d;
  wire                uSystolicPE_345_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_345_io_randW_d;
  wire       [14:0]   uSystolicPE_345_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_345_io_ofm_d;
  wire                uSystolicPE_346_io_mac_done_d;
  wire                uSystolicPE_346_io_enable_i_d;
  wire                uSystolicPE_346_io_clear_i_d;
  wire                uSystolicPE_346_io_enable_w_d;
  wire                uSystolicPE_346_io_clear_w_d;
  wire                uSystolicPE_346_io_enable_o_d;
  wire                uSystolicPE_346_io_clear_o_d;
  wire                uSystolicPE_346_io_ifm_sign_d;
  wire                uSystolicPE_346_io_ifm_dff_d;
  wire                uSystolicPE_346_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_346_io_randW_d;
  wire       [14:0]   uSystolicPE_346_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_346_io_ofm_d;
  wire                uSystolicPE_347_io_mac_done_d;
  wire                uSystolicPE_347_io_enable_i_d;
  wire                uSystolicPE_347_io_clear_i_d;
  wire                uSystolicPE_347_io_enable_w_d;
  wire                uSystolicPE_347_io_clear_w_d;
  wire                uSystolicPE_347_io_enable_o_d;
  wire                uSystolicPE_347_io_clear_o_d;
  wire                uSystolicPE_347_io_ifm_sign_d;
  wire                uSystolicPE_347_io_ifm_dff_d;
  wire                uSystolicPE_347_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_347_io_randW_d;
  wire       [14:0]   uSystolicPE_347_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_347_io_ofm_d;
  wire                uSystolicPE_348_io_mac_done_d;
  wire                uSystolicPE_348_io_enable_i_d;
  wire                uSystolicPE_348_io_clear_i_d;
  wire                uSystolicPE_348_io_enable_w_d;
  wire                uSystolicPE_348_io_clear_w_d;
  wire                uSystolicPE_348_io_enable_o_d;
  wire                uSystolicPE_348_io_clear_o_d;
  wire                uSystolicPE_348_io_ifm_sign_d;
  wire                uSystolicPE_348_io_ifm_dff_d;
  wire                uSystolicPE_348_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_348_io_randW_d;
  wire       [14:0]   uSystolicPE_348_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_348_io_ofm_d;
  wire                uSystolicPE_349_io_mac_done_d;
  wire                uSystolicPE_349_io_enable_i_d;
  wire                uSystolicPE_349_io_clear_i_d;
  wire                uSystolicPE_349_io_enable_w_d;
  wire                uSystolicPE_349_io_clear_w_d;
  wire                uSystolicPE_349_io_enable_o_d;
  wire                uSystolicPE_349_io_clear_o_d;
  wire                uSystolicPE_349_io_ifm_sign_d;
  wire                uSystolicPE_349_io_ifm_dff_d;
  wire                uSystolicPE_349_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_349_io_randW_d;
  wire       [14:0]   uSystolicPE_349_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_349_io_ofm_d;
  wire                uSystolicPE_350_io_mac_done_d;
  wire                uSystolicPE_350_io_enable_i_d;
  wire                uSystolicPE_350_io_clear_i_d;
  wire                uSystolicPE_350_io_enable_w_d;
  wire                uSystolicPE_350_io_clear_w_d;
  wire                uSystolicPE_350_io_enable_o_d;
  wire                uSystolicPE_350_io_clear_o_d;
  wire                uSystolicPE_350_io_ifm_sign_d;
  wire                uSystolicPE_350_io_ifm_dff_d;
  wire                uSystolicPE_350_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_350_io_randW_d;
  wire       [14:0]   uSystolicPE_350_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_350_io_ofm_d;
  wire                uSystolicPE_351_io_mac_done_d;
  wire                uSystolicPE_351_io_enable_i_d;
  wire                uSystolicPE_351_io_clear_i_d;
  wire                uSystolicPE_351_io_enable_w_d;
  wire                uSystolicPE_351_io_clear_w_d;
  wire                uSystolicPE_351_io_enable_o_d;
  wire                uSystolicPE_351_io_clear_o_d;
  wire                uSystolicPE_351_io_ifm_sign_d;
  wire                uSystolicPE_351_io_ifm_dff_d;
  wire                uSystolicPE_351_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_351_io_randW_d;
  wire       [14:0]   uSystolicPE_351_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_351_io_ofm_d;
  wire                uSystolicPE_352_io_mac_done_d;
  wire                uSystolicPE_352_io_enable_i_d;
  wire                uSystolicPE_352_io_clear_i_d;
  wire                uSystolicPE_352_io_enable_w_d;
  wire                uSystolicPE_352_io_clear_w_d;
  wire                uSystolicPE_352_io_enable_o_d;
  wire                uSystolicPE_352_io_clear_o_d;
  wire                uSystolicPE_352_io_ifm_sign_d;
  wire                uSystolicPE_352_io_ifm_dff_d;
  wire                uSystolicPE_352_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_352_io_randW_d;
  wire       [14:0]   uSystolicPE_352_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_352_io_ofm_d;
  wire                uSystolicPE_353_io_mac_done_d;
  wire                uSystolicPE_353_io_enable_i_d;
  wire                uSystolicPE_353_io_clear_i_d;
  wire                uSystolicPE_353_io_enable_w_d;
  wire                uSystolicPE_353_io_clear_w_d;
  wire                uSystolicPE_353_io_enable_o_d;
  wire                uSystolicPE_353_io_clear_o_d;
  wire                uSystolicPE_353_io_ifm_sign_d;
  wire                uSystolicPE_353_io_ifm_dff_d;
  wire                uSystolicPE_353_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_353_io_randW_d;
  wire       [14:0]   uSystolicPE_353_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_353_io_ofm_d;
  wire                uSystolicPE_354_io_mac_done_d;
  wire                uSystolicPE_354_io_enable_i_d;
  wire                uSystolicPE_354_io_clear_i_d;
  wire                uSystolicPE_354_io_enable_w_d;
  wire                uSystolicPE_354_io_clear_w_d;
  wire                uSystolicPE_354_io_enable_o_d;
  wire                uSystolicPE_354_io_clear_o_d;
  wire                uSystolicPE_354_io_ifm_sign_d;
  wire                uSystolicPE_354_io_ifm_dff_d;
  wire                uSystolicPE_354_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_354_io_randW_d;
  wire       [14:0]   uSystolicPE_354_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_354_io_ofm_d;
  wire                uSystolicPE_355_io_mac_done_d;
  wire                uSystolicPE_355_io_enable_i_d;
  wire                uSystolicPE_355_io_clear_i_d;
  wire                uSystolicPE_355_io_enable_w_d;
  wire                uSystolicPE_355_io_clear_w_d;
  wire                uSystolicPE_355_io_enable_o_d;
  wire                uSystolicPE_355_io_clear_o_d;
  wire                uSystolicPE_355_io_ifm_sign_d;
  wire                uSystolicPE_355_io_ifm_dff_d;
  wire                uSystolicPE_355_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_355_io_randW_d;
  wire       [14:0]   uSystolicPE_355_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_355_io_ofm_d;
  wire                uSystolicPE_356_io_mac_done_d;
  wire                uSystolicPE_356_io_enable_i_d;
  wire                uSystolicPE_356_io_clear_i_d;
  wire                uSystolicPE_356_io_enable_w_d;
  wire                uSystolicPE_356_io_clear_w_d;
  wire                uSystolicPE_356_io_enable_o_d;
  wire                uSystolicPE_356_io_clear_o_d;
  wire                uSystolicPE_356_io_ifm_sign_d;
  wire                uSystolicPE_356_io_ifm_dff_d;
  wire                uSystolicPE_356_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_356_io_randW_d;
  wire       [14:0]   uSystolicPE_356_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_356_io_ofm_d;
  wire                uSystolicPE_357_io_mac_done_d;
  wire                uSystolicPE_357_io_enable_i_d;
  wire                uSystolicPE_357_io_clear_i_d;
  wire                uSystolicPE_357_io_enable_w_d;
  wire                uSystolicPE_357_io_clear_w_d;
  wire                uSystolicPE_357_io_enable_o_d;
  wire                uSystolicPE_357_io_clear_o_d;
  wire                uSystolicPE_357_io_ifm_sign_d;
  wire                uSystolicPE_357_io_ifm_dff_d;
  wire                uSystolicPE_357_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_357_io_randW_d;
  wire       [14:0]   uSystolicPE_357_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_357_io_ofm_d;
  wire                uSystolicPE_358_io_mac_done_d;
  wire                uSystolicPE_358_io_enable_i_d;
  wire                uSystolicPE_358_io_clear_i_d;
  wire                uSystolicPE_358_io_enable_w_d;
  wire                uSystolicPE_358_io_clear_w_d;
  wire                uSystolicPE_358_io_enable_o_d;
  wire                uSystolicPE_358_io_clear_o_d;
  wire                uSystolicPE_358_io_ifm_sign_d;
  wire                uSystolicPE_358_io_ifm_dff_d;
  wire                uSystolicPE_358_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_358_io_randW_d;
  wire       [14:0]   uSystolicPE_358_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_358_io_ofm_d;
  wire                uSystolicPE_359_io_mac_done_d;
  wire                uSystolicPE_359_io_enable_i_d;
  wire                uSystolicPE_359_io_clear_i_d;
  wire                uSystolicPE_359_io_enable_w_d;
  wire                uSystolicPE_359_io_clear_w_d;
  wire                uSystolicPE_359_io_enable_o_d;
  wire                uSystolicPE_359_io_clear_o_d;
  wire                uSystolicPE_359_io_ifm_sign_d;
  wire                uSystolicPE_359_io_ifm_dff_d;
  wire                uSystolicPE_359_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_359_io_randW_d;
  wire       [14:0]   uSystolicPE_359_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_359_io_ofm_d;
  wire                uSystolicPEBorder_24_io_mac_done_d;
  wire                uSystolicPEBorder_24_io_enable_i_d;
  wire                uSystolicPEBorder_24_io_clear_i_d;
  wire                uSystolicPEBorder_24_io_enable_w_d;
  wire                uSystolicPEBorder_24_io_clear_w_d;
  wire                uSystolicPEBorder_24_io_enable_o_d;
  wire                uSystolicPEBorder_24_io_clear_o_d;
  wire                uSystolicPEBorder_24_io_ifm_sign_d;
  wire                uSystolicPEBorder_24_io_ifm_dff_d;
  wire                uSystolicPEBorder_24_io_wght_sign_d;
  wire       [14:0]   uSystolicPEBorder_24_io_randW_d;
  wire       [14:0]   uSystolicPEBorder_24_io_wght_abs_d;
  wire       [31:0]   uSystolicPEBorder_24_io_ofm_d;
  wire                uSystolicPE_360_io_mac_done_d;
  wire                uSystolicPE_360_io_enable_i_d;
  wire                uSystolicPE_360_io_clear_i_d;
  wire                uSystolicPE_360_io_enable_w_d;
  wire                uSystolicPE_360_io_clear_w_d;
  wire                uSystolicPE_360_io_enable_o_d;
  wire                uSystolicPE_360_io_clear_o_d;
  wire                uSystolicPE_360_io_ifm_sign_d;
  wire                uSystolicPE_360_io_ifm_dff_d;
  wire                uSystolicPE_360_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_360_io_randW_d;
  wire       [14:0]   uSystolicPE_360_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_360_io_ofm_d;
  wire                uSystolicPE_361_io_mac_done_d;
  wire                uSystolicPE_361_io_enable_i_d;
  wire                uSystolicPE_361_io_clear_i_d;
  wire                uSystolicPE_361_io_enable_w_d;
  wire                uSystolicPE_361_io_clear_w_d;
  wire                uSystolicPE_361_io_enable_o_d;
  wire                uSystolicPE_361_io_clear_o_d;
  wire                uSystolicPE_361_io_ifm_sign_d;
  wire                uSystolicPE_361_io_ifm_dff_d;
  wire                uSystolicPE_361_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_361_io_randW_d;
  wire       [14:0]   uSystolicPE_361_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_361_io_ofm_d;
  wire                uSystolicPE_362_io_mac_done_d;
  wire                uSystolicPE_362_io_enable_i_d;
  wire                uSystolicPE_362_io_clear_i_d;
  wire                uSystolicPE_362_io_enable_w_d;
  wire                uSystolicPE_362_io_clear_w_d;
  wire                uSystolicPE_362_io_enable_o_d;
  wire                uSystolicPE_362_io_clear_o_d;
  wire                uSystolicPE_362_io_ifm_sign_d;
  wire                uSystolicPE_362_io_ifm_dff_d;
  wire                uSystolicPE_362_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_362_io_randW_d;
  wire       [14:0]   uSystolicPE_362_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_362_io_ofm_d;
  wire                uSystolicPE_363_io_mac_done_d;
  wire                uSystolicPE_363_io_enable_i_d;
  wire                uSystolicPE_363_io_clear_i_d;
  wire                uSystolicPE_363_io_enable_w_d;
  wire                uSystolicPE_363_io_clear_w_d;
  wire                uSystolicPE_363_io_enable_o_d;
  wire                uSystolicPE_363_io_clear_o_d;
  wire                uSystolicPE_363_io_ifm_sign_d;
  wire                uSystolicPE_363_io_ifm_dff_d;
  wire                uSystolicPE_363_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_363_io_randW_d;
  wire       [14:0]   uSystolicPE_363_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_363_io_ofm_d;
  wire                uSystolicPE_364_io_mac_done_d;
  wire                uSystolicPE_364_io_enable_i_d;
  wire                uSystolicPE_364_io_clear_i_d;
  wire                uSystolicPE_364_io_enable_w_d;
  wire                uSystolicPE_364_io_clear_w_d;
  wire                uSystolicPE_364_io_enable_o_d;
  wire                uSystolicPE_364_io_clear_o_d;
  wire                uSystolicPE_364_io_ifm_sign_d;
  wire                uSystolicPE_364_io_ifm_dff_d;
  wire                uSystolicPE_364_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_364_io_randW_d;
  wire       [14:0]   uSystolicPE_364_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_364_io_ofm_d;
  wire                uSystolicPE_365_io_mac_done_d;
  wire                uSystolicPE_365_io_enable_i_d;
  wire                uSystolicPE_365_io_clear_i_d;
  wire                uSystolicPE_365_io_enable_w_d;
  wire                uSystolicPE_365_io_clear_w_d;
  wire                uSystolicPE_365_io_enable_o_d;
  wire                uSystolicPE_365_io_clear_o_d;
  wire                uSystolicPE_365_io_ifm_sign_d;
  wire                uSystolicPE_365_io_ifm_dff_d;
  wire                uSystolicPE_365_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_365_io_randW_d;
  wire       [14:0]   uSystolicPE_365_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_365_io_ofm_d;
  wire                uSystolicPE_366_io_mac_done_d;
  wire                uSystolicPE_366_io_enable_i_d;
  wire                uSystolicPE_366_io_clear_i_d;
  wire                uSystolicPE_366_io_enable_w_d;
  wire                uSystolicPE_366_io_clear_w_d;
  wire                uSystolicPE_366_io_enable_o_d;
  wire                uSystolicPE_366_io_clear_o_d;
  wire                uSystolicPE_366_io_ifm_sign_d;
  wire                uSystolicPE_366_io_ifm_dff_d;
  wire                uSystolicPE_366_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_366_io_randW_d;
  wire       [14:0]   uSystolicPE_366_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_366_io_ofm_d;
  wire                uSystolicPE_367_io_mac_done_d;
  wire                uSystolicPE_367_io_enable_i_d;
  wire                uSystolicPE_367_io_clear_i_d;
  wire                uSystolicPE_367_io_enable_w_d;
  wire                uSystolicPE_367_io_clear_w_d;
  wire                uSystolicPE_367_io_enable_o_d;
  wire                uSystolicPE_367_io_clear_o_d;
  wire                uSystolicPE_367_io_ifm_sign_d;
  wire                uSystolicPE_367_io_ifm_dff_d;
  wire                uSystolicPE_367_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_367_io_randW_d;
  wire       [14:0]   uSystolicPE_367_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_367_io_ofm_d;
  wire                uSystolicPE_368_io_mac_done_d;
  wire                uSystolicPE_368_io_enable_i_d;
  wire                uSystolicPE_368_io_clear_i_d;
  wire                uSystolicPE_368_io_enable_w_d;
  wire                uSystolicPE_368_io_clear_w_d;
  wire                uSystolicPE_368_io_enable_o_d;
  wire                uSystolicPE_368_io_clear_o_d;
  wire                uSystolicPE_368_io_ifm_sign_d;
  wire                uSystolicPE_368_io_ifm_dff_d;
  wire                uSystolicPE_368_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_368_io_randW_d;
  wire       [14:0]   uSystolicPE_368_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_368_io_ofm_d;
  wire                uSystolicPE_369_io_mac_done_d;
  wire                uSystolicPE_369_io_enable_i_d;
  wire                uSystolicPE_369_io_clear_i_d;
  wire                uSystolicPE_369_io_enable_w_d;
  wire                uSystolicPE_369_io_clear_w_d;
  wire                uSystolicPE_369_io_enable_o_d;
  wire                uSystolicPE_369_io_clear_o_d;
  wire                uSystolicPE_369_io_ifm_sign_d;
  wire                uSystolicPE_369_io_ifm_dff_d;
  wire                uSystolicPE_369_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_369_io_randW_d;
  wire       [14:0]   uSystolicPE_369_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_369_io_ofm_d;
  wire                uSystolicPE_370_io_mac_done_d;
  wire                uSystolicPE_370_io_enable_i_d;
  wire                uSystolicPE_370_io_clear_i_d;
  wire                uSystolicPE_370_io_enable_w_d;
  wire                uSystolicPE_370_io_clear_w_d;
  wire                uSystolicPE_370_io_enable_o_d;
  wire                uSystolicPE_370_io_clear_o_d;
  wire                uSystolicPE_370_io_ifm_sign_d;
  wire                uSystolicPE_370_io_ifm_dff_d;
  wire                uSystolicPE_370_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_370_io_randW_d;
  wire       [14:0]   uSystolicPE_370_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_370_io_ofm_d;
  wire                uSystolicPE_371_io_mac_done_d;
  wire                uSystolicPE_371_io_enable_i_d;
  wire                uSystolicPE_371_io_clear_i_d;
  wire                uSystolicPE_371_io_enable_w_d;
  wire                uSystolicPE_371_io_clear_w_d;
  wire                uSystolicPE_371_io_enable_o_d;
  wire                uSystolicPE_371_io_clear_o_d;
  wire                uSystolicPE_371_io_ifm_sign_d;
  wire                uSystolicPE_371_io_ifm_dff_d;
  wire                uSystolicPE_371_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_371_io_randW_d;
  wire       [14:0]   uSystolicPE_371_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_371_io_ofm_d;
  wire                uSystolicPE_372_io_mac_done_d;
  wire                uSystolicPE_372_io_enable_i_d;
  wire                uSystolicPE_372_io_clear_i_d;
  wire                uSystolicPE_372_io_enable_w_d;
  wire                uSystolicPE_372_io_clear_w_d;
  wire                uSystolicPE_372_io_enable_o_d;
  wire                uSystolicPE_372_io_clear_o_d;
  wire                uSystolicPE_372_io_ifm_sign_d;
  wire                uSystolicPE_372_io_ifm_dff_d;
  wire                uSystolicPE_372_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_372_io_randW_d;
  wire       [14:0]   uSystolicPE_372_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_372_io_ofm_d;
  wire                uSystolicPE_373_io_mac_done_d;
  wire                uSystolicPE_373_io_enable_i_d;
  wire                uSystolicPE_373_io_clear_i_d;
  wire                uSystolicPE_373_io_enable_w_d;
  wire                uSystolicPE_373_io_clear_w_d;
  wire                uSystolicPE_373_io_enable_o_d;
  wire                uSystolicPE_373_io_clear_o_d;
  wire                uSystolicPE_373_io_ifm_sign_d;
  wire                uSystolicPE_373_io_ifm_dff_d;
  wire                uSystolicPE_373_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_373_io_randW_d;
  wire       [14:0]   uSystolicPE_373_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_373_io_ofm_d;
  wire                uSystolicPE_374_io_mac_done_d;
  wire                uSystolicPE_374_io_enable_i_d;
  wire                uSystolicPE_374_io_clear_i_d;
  wire                uSystolicPE_374_io_enable_w_d;
  wire                uSystolicPE_374_io_clear_w_d;
  wire                uSystolicPE_374_io_enable_o_d;
  wire                uSystolicPE_374_io_clear_o_d;
  wire                uSystolicPE_374_io_ifm_sign_d;
  wire                uSystolicPE_374_io_ifm_dff_d;
  wire                uSystolicPE_374_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_374_io_randW_d;
  wire       [14:0]   uSystolicPE_374_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_374_io_ofm_d;
  wire                uSystolicPEBorder_25_io_mac_done_d;
  wire                uSystolicPEBorder_25_io_enable_i_d;
  wire                uSystolicPEBorder_25_io_clear_i_d;
  wire                uSystolicPEBorder_25_io_enable_w_d;
  wire                uSystolicPEBorder_25_io_clear_w_d;
  wire                uSystolicPEBorder_25_io_enable_o_d;
  wire                uSystolicPEBorder_25_io_clear_o_d;
  wire                uSystolicPEBorder_25_io_ifm_sign_d;
  wire                uSystolicPEBorder_25_io_ifm_dff_d;
  wire                uSystolicPEBorder_25_io_wght_sign_d;
  wire       [14:0]   uSystolicPEBorder_25_io_randW_d;
  wire       [14:0]   uSystolicPEBorder_25_io_wght_abs_d;
  wire       [31:0]   uSystolicPEBorder_25_io_ofm_d;
  wire                uSystolicPE_375_io_mac_done_d;
  wire                uSystolicPE_375_io_enable_i_d;
  wire                uSystolicPE_375_io_clear_i_d;
  wire                uSystolicPE_375_io_enable_w_d;
  wire                uSystolicPE_375_io_clear_w_d;
  wire                uSystolicPE_375_io_enable_o_d;
  wire                uSystolicPE_375_io_clear_o_d;
  wire                uSystolicPE_375_io_ifm_sign_d;
  wire                uSystolicPE_375_io_ifm_dff_d;
  wire                uSystolicPE_375_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_375_io_randW_d;
  wire       [14:0]   uSystolicPE_375_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_375_io_ofm_d;
  wire                uSystolicPE_376_io_mac_done_d;
  wire                uSystolicPE_376_io_enable_i_d;
  wire                uSystolicPE_376_io_clear_i_d;
  wire                uSystolicPE_376_io_enable_w_d;
  wire                uSystolicPE_376_io_clear_w_d;
  wire                uSystolicPE_376_io_enable_o_d;
  wire                uSystolicPE_376_io_clear_o_d;
  wire                uSystolicPE_376_io_ifm_sign_d;
  wire                uSystolicPE_376_io_ifm_dff_d;
  wire                uSystolicPE_376_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_376_io_randW_d;
  wire       [14:0]   uSystolicPE_376_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_376_io_ofm_d;
  wire                uSystolicPE_377_io_mac_done_d;
  wire                uSystolicPE_377_io_enable_i_d;
  wire                uSystolicPE_377_io_clear_i_d;
  wire                uSystolicPE_377_io_enable_w_d;
  wire                uSystolicPE_377_io_clear_w_d;
  wire                uSystolicPE_377_io_enable_o_d;
  wire                uSystolicPE_377_io_clear_o_d;
  wire                uSystolicPE_377_io_ifm_sign_d;
  wire                uSystolicPE_377_io_ifm_dff_d;
  wire                uSystolicPE_377_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_377_io_randW_d;
  wire       [14:0]   uSystolicPE_377_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_377_io_ofm_d;
  wire                uSystolicPE_378_io_mac_done_d;
  wire                uSystolicPE_378_io_enable_i_d;
  wire                uSystolicPE_378_io_clear_i_d;
  wire                uSystolicPE_378_io_enable_w_d;
  wire                uSystolicPE_378_io_clear_w_d;
  wire                uSystolicPE_378_io_enable_o_d;
  wire                uSystolicPE_378_io_clear_o_d;
  wire                uSystolicPE_378_io_ifm_sign_d;
  wire                uSystolicPE_378_io_ifm_dff_d;
  wire                uSystolicPE_378_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_378_io_randW_d;
  wire       [14:0]   uSystolicPE_378_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_378_io_ofm_d;
  wire                uSystolicPE_379_io_mac_done_d;
  wire                uSystolicPE_379_io_enable_i_d;
  wire                uSystolicPE_379_io_clear_i_d;
  wire                uSystolicPE_379_io_enable_w_d;
  wire                uSystolicPE_379_io_clear_w_d;
  wire                uSystolicPE_379_io_enable_o_d;
  wire                uSystolicPE_379_io_clear_o_d;
  wire                uSystolicPE_379_io_ifm_sign_d;
  wire                uSystolicPE_379_io_ifm_dff_d;
  wire                uSystolicPE_379_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_379_io_randW_d;
  wire       [14:0]   uSystolicPE_379_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_379_io_ofm_d;
  wire                uSystolicPE_380_io_mac_done_d;
  wire                uSystolicPE_380_io_enable_i_d;
  wire                uSystolicPE_380_io_clear_i_d;
  wire                uSystolicPE_380_io_enable_w_d;
  wire                uSystolicPE_380_io_clear_w_d;
  wire                uSystolicPE_380_io_enable_o_d;
  wire                uSystolicPE_380_io_clear_o_d;
  wire                uSystolicPE_380_io_ifm_sign_d;
  wire                uSystolicPE_380_io_ifm_dff_d;
  wire                uSystolicPE_380_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_380_io_randW_d;
  wire       [14:0]   uSystolicPE_380_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_380_io_ofm_d;
  wire                uSystolicPE_381_io_mac_done_d;
  wire                uSystolicPE_381_io_enable_i_d;
  wire                uSystolicPE_381_io_clear_i_d;
  wire                uSystolicPE_381_io_enable_w_d;
  wire                uSystolicPE_381_io_clear_w_d;
  wire                uSystolicPE_381_io_enable_o_d;
  wire                uSystolicPE_381_io_clear_o_d;
  wire                uSystolicPE_381_io_ifm_sign_d;
  wire                uSystolicPE_381_io_ifm_dff_d;
  wire                uSystolicPE_381_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_381_io_randW_d;
  wire       [14:0]   uSystolicPE_381_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_381_io_ofm_d;
  wire                uSystolicPE_382_io_mac_done_d;
  wire                uSystolicPE_382_io_enable_i_d;
  wire                uSystolicPE_382_io_clear_i_d;
  wire                uSystolicPE_382_io_enable_w_d;
  wire                uSystolicPE_382_io_clear_w_d;
  wire                uSystolicPE_382_io_enable_o_d;
  wire                uSystolicPE_382_io_clear_o_d;
  wire                uSystolicPE_382_io_ifm_sign_d;
  wire                uSystolicPE_382_io_ifm_dff_d;
  wire                uSystolicPE_382_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_382_io_randW_d;
  wire       [14:0]   uSystolicPE_382_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_382_io_ofm_d;
  wire                uSystolicPE_383_io_mac_done_d;
  wire                uSystolicPE_383_io_enable_i_d;
  wire                uSystolicPE_383_io_clear_i_d;
  wire                uSystolicPE_383_io_enable_w_d;
  wire                uSystolicPE_383_io_clear_w_d;
  wire                uSystolicPE_383_io_enable_o_d;
  wire                uSystolicPE_383_io_clear_o_d;
  wire                uSystolicPE_383_io_ifm_sign_d;
  wire                uSystolicPE_383_io_ifm_dff_d;
  wire                uSystolicPE_383_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_383_io_randW_d;
  wire       [14:0]   uSystolicPE_383_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_383_io_ofm_d;
  wire                uSystolicPE_384_io_mac_done_d;
  wire                uSystolicPE_384_io_enable_i_d;
  wire                uSystolicPE_384_io_clear_i_d;
  wire                uSystolicPE_384_io_enable_w_d;
  wire                uSystolicPE_384_io_clear_w_d;
  wire                uSystolicPE_384_io_enable_o_d;
  wire                uSystolicPE_384_io_clear_o_d;
  wire                uSystolicPE_384_io_ifm_sign_d;
  wire                uSystolicPE_384_io_ifm_dff_d;
  wire                uSystolicPE_384_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_384_io_randW_d;
  wire       [14:0]   uSystolicPE_384_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_384_io_ofm_d;
  wire                uSystolicPE_385_io_mac_done_d;
  wire                uSystolicPE_385_io_enable_i_d;
  wire                uSystolicPE_385_io_clear_i_d;
  wire                uSystolicPE_385_io_enable_w_d;
  wire                uSystolicPE_385_io_clear_w_d;
  wire                uSystolicPE_385_io_enable_o_d;
  wire                uSystolicPE_385_io_clear_o_d;
  wire                uSystolicPE_385_io_ifm_sign_d;
  wire                uSystolicPE_385_io_ifm_dff_d;
  wire                uSystolicPE_385_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_385_io_randW_d;
  wire       [14:0]   uSystolicPE_385_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_385_io_ofm_d;
  wire                uSystolicPE_386_io_mac_done_d;
  wire                uSystolicPE_386_io_enable_i_d;
  wire                uSystolicPE_386_io_clear_i_d;
  wire                uSystolicPE_386_io_enable_w_d;
  wire                uSystolicPE_386_io_clear_w_d;
  wire                uSystolicPE_386_io_enable_o_d;
  wire                uSystolicPE_386_io_clear_o_d;
  wire                uSystolicPE_386_io_ifm_sign_d;
  wire                uSystolicPE_386_io_ifm_dff_d;
  wire                uSystolicPE_386_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_386_io_randW_d;
  wire       [14:0]   uSystolicPE_386_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_386_io_ofm_d;
  wire                uSystolicPE_387_io_mac_done_d;
  wire                uSystolicPE_387_io_enable_i_d;
  wire                uSystolicPE_387_io_clear_i_d;
  wire                uSystolicPE_387_io_enable_w_d;
  wire                uSystolicPE_387_io_clear_w_d;
  wire                uSystolicPE_387_io_enable_o_d;
  wire                uSystolicPE_387_io_clear_o_d;
  wire                uSystolicPE_387_io_ifm_sign_d;
  wire                uSystolicPE_387_io_ifm_dff_d;
  wire                uSystolicPE_387_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_387_io_randW_d;
  wire       [14:0]   uSystolicPE_387_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_387_io_ofm_d;
  wire                uSystolicPE_388_io_mac_done_d;
  wire                uSystolicPE_388_io_enable_i_d;
  wire                uSystolicPE_388_io_clear_i_d;
  wire                uSystolicPE_388_io_enable_w_d;
  wire                uSystolicPE_388_io_clear_w_d;
  wire                uSystolicPE_388_io_enable_o_d;
  wire                uSystolicPE_388_io_clear_o_d;
  wire                uSystolicPE_388_io_ifm_sign_d;
  wire                uSystolicPE_388_io_ifm_dff_d;
  wire                uSystolicPE_388_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_388_io_randW_d;
  wire       [14:0]   uSystolicPE_388_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_388_io_ofm_d;
  wire                uSystolicPE_389_io_mac_done_d;
  wire                uSystolicPE_389_io_enable_i_d;
  wire                uSystolicPE_389_io_clear_i_d;
  wire                uSystolicPE_389_io_enable_w_d;
  wire                uSystolicPE_389_io_clear_w_d;
  wire                uSystolicPE_389_io_enable_o_d;
  wire                uSystolicPE_389_io_clear_o_d;
  wire                uSystolicPE_389_io_ifm_sign_d;
  wire                uSystolicPE_389_io_ifm_dff_d;
  wire                uSystolicPE_389_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_389_io_randW_d;
  wire       [14:0]   uSystolicPE_389_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_389_io_ofm_d;
  wire                uSystolicPEBorder_26_io_mac_done_d;
  wire                uSystolicPEBorder_26_io_enable_i_d;
  wire                uSystolicPEBorder_26_io_clear_i_d;
  wire                uSystolicPEBorder_26_io_enable_w_d;
  wire                uSystolicPEBorder_26_io_clear_w_d;
  wire                uSystolicPEBorder_26_io_enable_o_d;
  wire                uSystolicPEBorder_26_io_clear_o_d;
  wire                uSystolicPEBorder_26_io_ifm_sign_d;
  wire                uSystolicPEBorder_26_io_ifm_dff_d;
  wire                uSystolicPEBorder_26_io_wght_sign_d;
  wire       [14:0]   uSystolicPEBorder_26_io_randW_d;
  wire       [14:0]   uSystolicPEBorder_26_io_wght_abs_d;
  wire       [31:0]   uSystolicPEBorder_26_io_ofm_d;
  wire                uSystolicPE_390_io_mac_done_d;
  wire                uSystolicPE_390_io_enable_i_d;
  wire                uSystolicPE_390_io_clear_i_d;
  wire                uSystolicPE_390_io_enable_w_d;
  wire                uSystolicPE_390_io_clear_w_d;
  wire                uSystolicPE_390_io_enable_o_d;
  wire                uSystolicPE_390_io_clear_o_d;
  wire                uSystolicPE_390_io_ifm_sign_d;
  wire                uSystolicPE_390_io_ifm_dff_d;
  wire                uSystolicPE_390_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_390_io_randW_d;
  wire       [14:0]   uSystolicPE_390_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_390_io_ofm_d;
  wire                uSystolicPE_391_io_mac_done_d;
  wire                uSystolicPE_391_io_enable_i_d;
  wire                uSystolicPE_391_io_clear_i_d;
  wire                uSystolicPE_391_io_enable_w_d;
  wire                uSystolicPE_391_io_clear_w_d;
  wire                uSystolicPE_391_io_enable_o_d;
  wire                uSystolicPE_391_io_clear_o_d;
  wire                uSystolicPE_391_io_ifm_sign_d;
  wire                uSystolicPE_391_io_ifm_dff_d;
  wire                uSystolicPE_391_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_391_io_randW_d;
  wire       [14:0]   uSystolicPE_391_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_391_io_ofm_d;
  wire                uSystolicPE_392_io_mac_done_d;
  wire                uSystolicPE_392_io_enable_i_d;
  wire                uSystolicPE_392_io_clear_i_d;
  wire                uSystolicPE_392_io_enable_w_d;
  wire                uSystolicPE_392_io_clear_w_d;
  wire                uSystolicPE_392_io_enable_o_d;
  wire                uSystolicPE_392_io_clear_o_d;
  wire                uSystolicPE_392_io_ifm_sign_d;
  wire                uSystolicPE_392_io_ifm_dff_d;
  wire                uSystolicPE_392_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_392_io_randW_d;
  wire       [14:0]   uSystolicPE_392_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_392_io_ofm_d;
  wire                uSystolicPE_393_io_mac_done_d;
  wire                uSystolicPE_393_io_enable_i_d;
  wire                uSystolicPE_393_io_clear_i_d;
  wire                uSystolicPE_393_io_enable_w_d;
  wire                uSystolicPE_393_io_clear_w_d;
  wire                uSystolicPE_393_io_enable_o_d;
  wire                uSystolicPE_393_io_clear_o_d;
  wire                uSystolicPE_393_io_ifm_sign_d;
  wire                uSystolicPE_393_io_ifm_dff_d;
  wire                uSystolicPE_393_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_393_io_randW_d;
  wire       [14:0]   uSystolicPE_393_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_393_io_ofm_d;
  wire                uSystolicPE_394_io_mac_done_d;
  wire                uSystolicPE_394_io_enable_i_d;
  wire                uSystolicPE_394_io_clear_i_d;
  wire                uSystolicPE_394_io_enable_w_d;
  wire                uSystolicPE_394_io_clear_w_d;
  wire                uSystolicPE_394_io_enable_o_d;
  wire                uSystolicPE_394_io_clear_o_d;
  wire                uSystolicPE_394_io_ifm_sign_d;
  wire                uSystolicPE_394_io_ifm_dff_d;
  wire                uSystolicPE_394_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_394_io_randW_d;
  wire       [14:0]   uSystolicPE_394_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_394_io_ofm_d;
  wire                uSystolicPE_395_io_mac_done_d;
  wire                uSystolicPE_395_io_enable_i_d;
  wire                uSystolicPE_395_io_clear_i_d;
  wire                uSystolicPE_395_io_enable_w_d;
  wire                uSystolicPE_395_io_clear_w_d;
  wire                uSystolicPE_395_io_enable_o_d;
  wire                uSystolicPE_395_io_clear_o_d;
  wire                uSystolicPE_395_io_ifm_sign_d;
  wire                uSystolicPE_395_io_ifm_dff_d;
  wire                uSystolicPE_395_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_395_io_randW_d;
  wire       [14:0]   uSystolicPE_395_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_395_io_ofm_d;
  wire                uSystolicPE_396_io_mac_done_d;
  wire                uSystolicPE_396_io_enable_i_d;
  wire                uSystolicPE_396_io_clear_i_d;
  wire                uSystolicPE_396_io_enable_w_d;
  wire                uSystolicPE_396_io_clear_w_d;
  wire                uSystolicPE_396_io_enable_o_d;
  wire                uSystolicPE_396_io_clear_o_d;
  wire                uSystolicPE_396_io_ifm_sign_d;
  wire                uSystolicPE_396_io_ifm_dff_d;
  wire                uSystolicPE_396_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_396_io_randW_d;
  wire       [14:0]   uSystolicPE_396_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_396_io_ofm_d;
  wire                uSystolicPE_397_io_mac_done_d;
  wire                uSystolicPE_397_io_enable_i_d;
  wire                uSystolicPE_397_io_clear_i_d;
  wire                uSystolicPE_397_io_enable_w_d;
  wire                uSystolicPE_397_io_clear_w_d;
  wire                uSystolicPE_397_io_enable_o_d;
  wire                uSystolicPE_397_io_clear_o_d;
  wire                uSystolicPE_397_io_ifm_sign_d;
  wire                uSystolicPE_397_io_ifm_dff_d;
  wire                uSystolicPE_397_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_397_io_randW_d;
  wire       [14:0]   uSystolicPE_397_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_397_io_ofm_d;
  wire                uSystolicPE_398_io_mac_done_d;
  wire                uSystolicPE_398_io_enable_i_d;
  wire                uSystolicPE_398_io_clear_i_d;
  wire                uSystolicPE_398_io_enable_w_d;
  wire                uSystolicPE_398_io_clear_w_d;
  wire                uSystolicPE_398_io_enable_o_d;
  wire                uSystolicPE_398_io_clear_o_d;
  wire                uSystolicPE_398_io_ifm_sign_d;
  wire                uSystolicPE_398_io_ifm_dff_d;
  wire                uSystolicPE_398_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_398_io_randW_d;
  wire       [14:0]   uSystolicPE_398_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_398_io_ofm_d;
  wire                uSystolicPE_399_io_mac_done_d;
  wire                uSystolicPE_399_io_enable_i_d;
  wire                uSystolicPE_399_io_clear_i_d;
  wire                uSystolicPE_399_io_enable_w_d;
  wire                uSystolicPE_399_io_clear_w_d;
  wire                uSystolicPE_399_io_enable_o_d;
  wire                uSystolicPE_399_io_clear_o_d;
  wire                uSystolicPE_399_io_ifm_sign_d;
  wire                uSystolicPE_399_io_ifm_dff_d;
  wire                uSystolicPE_399_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_399_io_randW_d;
  wire       [14:0]   uSystolicPE_399_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_399_io_ofm_d;
  wire                uSystolicPE_400_io_mac_done_d;
  wire                uSystolicPE_400_io_enable_i_d;
  wire                uSystolicPE_400_io_clear_i_d;
  wire                uSystolicPE_400_io_enable_w_d;
  wire                uSystolicPE_400_io_clear_w_d;
  wire                uSystolicPE_400_io_enable_o_d;
  wire                uSystolicPE_400_io_clear_o_d;
  wire                uSystolicPE_400_io_ifm_sign_d;
  wire                uSystolicPE_400_io_ifm_dff_d;
  wire                uSystolicPE_400_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_400_io_randW_d;
  wire       [14:0]   uSystolicPE_400_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_400_io_ofm_d;
  wire                uSystolicPE_401_io_mac_done_d;
  wire                uSystolicPE_401_io_enable_i_d;
  wire                uSystolicPE_401_io_clear_i_d;
  wire                uSystolicPE_401_io_enable_w_d;
  wire                uSystolicPE_401_io_clear_w_d;
  wire                uSystolicPE_401_io_enable_o_d;
  wire                uSystolicPE_401_io_clear_o_d;
  wire                uSystolicPE_401_io_ifm_sign_d;
  wire                uSystolicPE_401_io_ifm_dff_d;
  wire                uSystolicPE_401_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_401_io_randW_d;
  wire       [14:0]   uSystolicPE_401_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_401_io_ofm_d;
  wire                uSystolicPE_402_io_mac_done_d;
  wire                uSystolicPE_402_io_enable_i_d;
  wire                uSystolicPE_402_io_clear_i_d;
  wire                uSystolicPE_402_io_enable_w_d;
  wire                uSystolicPE_402_io_clear_w_d;
  wire                uSystolicPE_402_io_enable_o_d;
  wire                uSystolicPE_402_io_clear_o_d;
  wire                uSystolicPE_402_io_ifm_sign_d;
  wire                uSystolicPE_402_io_ifm_dff_d;
  wire                uSystolicPE_402_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_402_io_randW_d;
  wire       [14:0]   uSystolicPE_402_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_402_io_ofm_d;
  wire                uSystolicPE_403_io_mac_done_d;
  wire                uSystolicPE_403_io_enable_i_d;
  wire                uSystolicPE_403_io_clear_i_d;
  wire                uSystolicPE_403_io_enable_w_d;
  wire                uSystolicPE_403_io_clear_w_d;
  wire                uSystolicPE_403_io_enable_o_d;
  wire                uSystolicPE_403_io_clear_o_d;
  wire                uSystolicPE_403_io_ifm_sign_d;
  wire                uSystolicPE_403_io_ifm_dff_d;
  wire                uSystolicPE_403_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_403_io_randW_d;
  wire       [14:0]   uSystolicPE_403_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_403_io_ofm_d;
  wire                uSystolicPE_404_io_mac_done_d;
  wire                uSystolicPE_404_io_enable_i_d;
  wire                uSystolicPE_404_io_clear_i_d;
  wire                uSystolicPE_404_io_enable_w_d;
  wire                uSystolicPE_404_io_clear_w_d;
  wire                uSystolicPE_404_io_enable_o_d;
  wire                uSystolicPE_404_io_clear_o_d;
  wire                uSystolicPE_404_io_ifm_sign_d;
  wire                uSystolicPE_404_io_ifm_dff_d;
  wire                uSystolicPE_404_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_404_io_randW_d;
  wire       [14:0]   uSystolicPE_404_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_404_io_ofm_d;
  wire                uSystolicPEBorder_27_io_mac_done_d;
  wire                uSystolicPEBorder_27_io_enable_i_d;
  wire                uSystolicPEBorder_27_io_clear_i_d;
  wire                uSystolicPEBorder_27_io_enable_w_d;
  wire                uSystolicPEBorder_27_io_clear_w_d;
  wire                uSystolicPEBorder_27_io_enable_o_d;
  wire                uSystolicPEBorder_27_io_clear_o_d;
  wire                uSystolicPEBorder_27_io_ifm_sign_d;
  wire                uSystolicPEBorder_27_io_ifm_dff_d;
  wire                uSystolicPEBorder_27_io_wght_sign_d;
  wire       [14:0]   uSystolicPEBorder_27_io_randW_d;
  wire       [14:0]   uSystolicPEBorder_27_io_wght_abs_d;
  wire       [31:0]   uSystolicPEBorder_27_io_ofm_d;
  wire                uSystolicPE_405_io_mac_done_d;
  wire                uSystolicPE_405_io_enable_i_d;
  wire                uSystolicPE_405_io_clear_i_d;
  wire                uSystolicPE_405_io_enable_w_d;
  wire                uSystolicPE_405_io_clear_w_d;
  wire                uSystolicPE_405_io_enable_o_d;
  wire                uSystolicPE_405_io_clear_o_d;
  wire                uSystolicPE_405_io_ifm_sign_d;
  wire                uSystolicPE_405_io_ifm_dff_d;
  wire                uSystolicPE_405_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_405_io_randW_d;
  wire       [14:0]   uSystolicPE_405_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_405_io_ofm_d;
  wire                uSystolicPE_406_io_mac_done_d;
  wire                uSystolicPE_406_io_enable_i_d;
  wire                uSystolicPE_406_io_clear_i_d;
  wire                uSystolicPE_406_io_enable_w_d;
  wire                uSystolicPE_406_io_clear_w_d;
  wire                uSystolicPE_406_io_enable_o_d;
  wire                uSystolicPE_406_io_clear_o_d;
  wire                uSystolicPE_406_io_ifm_sign_d;
  wire                uSystolicPE_406_io_ifm_dff_d;
  wire                uSystolicPE_406_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_406_io_randW_d;
  wire       [14:0]   uSystolicPE_406_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_406_io_ofm_d;
  wire                uSystolicPE_407_io_mac_done_d;
  wire                uSystolicPE_407_io_enable_i_d;
  wire                uSystolicPE_407_io_clear_i_d;
  wire                uSystolicPE_407_io_enable_w_d;
  wire                uSystolicPE_407_io_clear_w_d;
  wire                uSystolicPE_407_io_enable_o_d;
  wire                uSystolicPE_407_io_clear_o_d;
  wire                uSystolicPE_407_io_ifm_sign_d;
  wire                uSystolicPE_407_io_ifm_dff_d;
  wire                uSystolicPE_407_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_407_io_randW_d;
  wire       [14:0]   uSystolicPE_407_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_407_io_ofm_d;
  wire                uSystolicPE_408_io_mac_done_d;
  wire                uSystolicPE_408_io_enable_i_d;
  wire                uSystolicPE_408_io_clear_i_d;
  wire                uSystolicPE_408_io_enable_w_d;
  wire                uSystolicPE_408_io_clear_w_d;
  wire                uSystolicPE_408_io_enable_o_d;
  wire                uSystolicPE_408_io_clear_o_d;
  wire                uSystolicPE_408_io_ifm_sign_d;
  wire                uSystolicPE_408_io_ifm_dff_d;
  wire                uSystolicPE_408_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_408_io_randW_d;
  wire       [14:0]   uSystolicPE_408_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_408_io_ofm_d;
  wire                uSystolicPE_409_io_mac_done_d;
  wire                uSystolicPE_409_io_enable_i_d;
  wire                uSystolicPE_409_io_clear_i_d;
  wire                uSystolicPE_409_io_enable_w_d;
  wire                uSystolicPE_409_io_clear_w_d;
  wire                uSystolicPE_409_io_enable_o_d;
  wire                uSystolicPE_409_io_clear_o_d;
  wire                uSystolicPE_409_io_ifm_sign_d;
  wire                uSystolicPE_409_io_ifm_dff_d;
  wire                uSystolicPE_409_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_409_io_randW_d;
  wire       [14:0]   uSystolicPE_409_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_409_io_ofm_d;
  wire                uSystolicPE_410_io_mac_done_d;
  wire                uSystolicPE_410_io_enable_i_d;
  wire                uSystolicPE_410_io_clear_i_d;
  wire                uSystolicPE_410_io_enable_w_d;
  wire                uSystolicPE_410_io_clear_w_d;
  wire                uSystolicPE_410_io_enable_o_d;
  wire                uSystolicPE_410_io_clear_o_d;
  wire                uSystolicPE_410_io_ifm_sign_d;
  wire                uSystolicPE_410_io_ifm_dff_d;
  wire                uSystolicPE_410_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_410_io_randW_d;
  wire       [14:0]   uSystolicPE_410_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_410_io_ofm_d;
  wire                uSystolicPE_411_io_mac_done_d;
  wire                uSystolicPE_411_io_enable_i_d;
  wire                uSystolicPE_411_io_clear_i_d;
  wire                uSystolicPE_411_io_enable_w_d;
  wire                uSystolicPE_411_io_clear_w_d;
  wire                uSystolicPE_411_io_enable_o_d;
  wire                uSystolicPE_411_io_clear_o_d;
  wire                uSystolicPE_411_io_ifm_sign_d;
  wire                uSystolicPE_411_io_ifm_dff_d;
  wire                uSystolicPE_411_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_411_io_randW_d;
  wire       [14:0]   uSystolicPE_411_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_411_io_ofm_d;
  wire                uSystolicPE_412_io_mac_done_d;
  wire                uSystolicPE_412_io_enable_i_d;
  wire                uSystolicPE_412_io_clear_i_d;
  wire                uSystolicPE_412_io_enable_w_d;
  wire                uSystolicPE_412_io_clear_w_d;
  wire                uSystolicPE_412_io_enable_o_d;
  wire                uSystolicPE_412_io_clear_o_d;
  wire                uSystolicPE_412_io_ifm_sign_d;
  wire                uSystolicPE_412_io_ifm_dff_d;
  wire                uSystolicPE_412_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_412_io_randW_d;
  wire       [14:0]   uSystolicPE_412_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_412_io_ofm_d;
  wire                uSystolicPE_413_io_mac_done_d;
  wire                uSystolicPE_413_io_enable_i_d;
  wire                uSystolicPE_413_io_clear_i_d;
  wire                uSystolicPE_413_io_enable_w_d;
  wire                uSystolicPE_413_io_clear_w_d;
  wire                uSystolicPE_413_io_enable_o_d;
  wire                uSystolicPE_413_io_clear_o_d;
  wire                uSystolicPE_413_io_ifm_sign_d;
  wire                uSystolicPE_413_io_ifm_dff_d;
  wire                uSystolicPE_413_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_413_io_randW_d;
  wire       [14:0]   uSystolicPE_413_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_413_io_ofm_d;
  wire                uSystolicPE_414_io_mac_done_d;
  wire                uSystolicPE_414_io_enable_i_d;
  wire                uSystolicPE_414_io_clear_i_d;
  wire                uSystolicPE_414_io_enable_w_d;
  wire                uSystolicPE_414_io_clear_w_d;
  wire                uSystolicPE_414_io_enable_o_d;
  wire                uSystolicPE_414_io_clear_o_d;
  wire                uSystolicPE_414_io_ifm_sign_d;
  wire                uSystolicPE_414_io_ifm_dff_d;
  wire                uSystolicPE_414_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_414_io_randW_d;
  wire       [14:0]   uSystolicPE_414_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_414_io_ofm_d;
  wire                uSystolicPE_415_io_mac_done_d;
  wire                uSystolicPE_415_io_enable_i_d;
  wire                uSystolicPE_415_io_clear_i_d;
  wire                uSystolicPE_415_io_enable_w_d;
  wire                uSystolicPE_415_io_clear_w_d;
  wire                uSystolicPE_415_io_enable_o_d;
  wire                uSystolicPE_415_io_clear_o_d;
  wire                uSystolicPE_415_io_ifm_sign_d;
  wire                uSystolicPE_415_io_ifm_dff_d;
  wire                uSystolicPE_415_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_415_io_randW_d;
  wire       [14:0]   uSystolicPE_415_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_415_io_ofm_d;
  wire                uSystolicPE_416_io_mac_done_d;
  wire                uSystolicPE_416_io_enable_i_d;
  wire                uSystolicPE_416_io_clear_i_d;
  wire                uSystolicPE_416_io_enable_w_d;
  wire                uSystolicPE_416_io_clear_w_d;
  wire                uSystolicPE_416_io_enable_o_d;
  wire                uSystolicPE_416_io_clear_o_d;
  wire                uSystolicPE_416_io_ifm_sign_d;
  wire                uSystolicPE_416_io_ifm_dff_d;
  wire                uSystolicPE_416_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_416_io_randW_d;
  wire       [14:0]   uSystolicPE_416_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_416_io_ofm_d;
  wire                uSystolicPE_417_io_mac_done_d;
  wire                uSystolicPE_417_io_enable_i_d;
  wire                uSystolicPE_417_io_clear_i_d;
  wire                uSystolicPE_417_io_enable_w_d;
  wire                uSystolicPE_417_io_clear_w_d;
  wire                uSystolicPE_417_io_enable_o_d;
  wire                uSystolicPE_417_io_clear_o_d;
  wire                uSystolicPE_417_io_ifm_sign_d;
  wire                uSystolicPE_417_io_ifm_dff_d;
  wire                uSystolicPE_417_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_417_io_randW_d;
  wire       [14:0]   uSystolicPE_417_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_417_io_ofm_d;
  wire                uSystolicPE_418_io_mac_done_d;
  wire                uSystolicPE_418_io_enable_i_d;
  wire                uSystolicPE_418_io_clear_i_d;
  wire                uSystolicPE_418_io_enable_w_d;
  wire                uSystolicPE_418_io_clear_w_d;
  wire                uSystolicPE_418_io_enable_o_d;
  wire                uSystolicPE_418_io_clear_o_d;
  wire                uSystolicPE_418_io_ifm_sign_d;
  wire                uSystolicPE_418_io_ifm_dff_d;
  wire                uSystolicPE_418_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_418_io_randW_d;
  wire       [14:0]   uSystolicPE_418_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_418_io_ofm_d;
  wire                uSystolicPE_419_io_mac_done_d;
  wire                uSystolicPE_419_io_enable_i_d;
  wire                uSystolicPE_419_io_clear_i_d;
  wire                uSystolicPE_419_io_enable_w_d;
  wire                uSystolicPE_419_io_clear_w_d;
  wire                uSystolicPE_419_io_enable_o_d;
  wire                uSystolicPE_419_io_clear_o_d;
  wire                uSystolicPE_419_io_ifm_sign_d;
  wire                uSystolicPE_419_io_ifm_dff_d;
  wire                uSystolicPE_419_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_419_io_randW_d;
  wire       [14:0]   uSystolicPE_419_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_419_io_ofm_d;
  wire                uSystolicPEBorder_28_io_mac_done_d;
  wire                uSystolicPEBorder_28_io_enable_i_d;
  wire                uSystolicPEBorder_28_io_clear_i_d;
  wire                uSystolicPEBorder_28_io_enable_w_d;
  wire                uSystolicPEBorder_28_io_clear_w_d;
  wire                uSystolicPEBorder_28_io_enable_o_d;
  wire                uSystolicPEBorder_28_io_clear_o_d;
  wire                uSystolicPEBorder_28_io_ifm_sign_d;
  wire                uSystolicPEBorder_28_io_ifm_dff_d;
  wire                uSystolicPEBorder_28_io_wght_sign_d;
  wire       [14:0]   uSystolicPEBorder_28_io_randW_d;
  wire       [14:0]   uSystolicPEBorder_28_io_wght_abs_d;
  wire       [31:0]   uSystolicPEBorder_28_io_ofm_d;
  wire                uSystolicPE_420_io_mac_done_d;
  wire                uSystolicPE_420_io_enable_i_d;
  wire                uSystolicPE_420_io_clear_i_d;
  wire                uSystolicPE_420_io_enable_w_d;
  wire                uSystolicPE_420_io_clear_w_d;
  wire                uSystolicPE_420_io_enable_o_d;
  wire                uSystolicPE_420_io_clear_o_d;
  wire                uSystolicPE_420_io_ifm_sign_d;
  wire                uSystolicPE_420_io_ifm_dff_d;
  wire                uSystolicPE_420_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_420_io_randW_d;
  wire       [14:0]   uSystolicPE_420_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_420_io_ofm_d;
  wire                uSystolicPE_421_io_mac_done_d;
  wire                uSystolicPE_421_io_enable_i_d;
  wire                uSystolicPE_421_io_clear_i_d;
  wire                uSystolicPE_421_io_enable_w_d;
  wire                uSystolicPE_421_io_clear_w_d;
  wire                uSystolicPE_421_io_enable_o_d;
  wire                uSystolicPE_421_io_clear_o_d;
  wire                uSystolicPE_421_io_ifm_sign_d;
  wire                uSystolicPE_421_io_ifm_dff_d;
  wire                uSystolicPE_421_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_421_io_randW_d;
  wire       [14:0]   uSystolicPE_421_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_421_io_ofm_d;
  wire                uSystolicPE_422_io_mac_done_d;
  wire                uSystolicPE_422_io_enable_i_d;
  wire                uSystolicPE_422_io_clear_i_d;
  wire                uSystolicPE_422_io_enable_w_d;
  wire                uSystolicPE_422_io_clear_w_d;
  wire                uSystolicPE_422_io_enable_o_d;
  wire                uSystolicPE_422_io_clear_o_d;
  wire                uSystolicPE_422_io_ifm_sign_d;
  wire                uSystolicPE_422_io_ifm_dff_d;
  wire                uSystolicPE_422_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_422_io_randW_d;
  wire       [14:0]   uSystolicPE_422_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_422_io_ofm_d;
  wire                uSystolicPE_423_io_mac_done_d;
  wire                uSystolicPE_423_io_enable_i_d;
  wire                uSystolicPE_423_io_clear_i_d;
  wire                uSystolicPE_423_io_enable_w_d;
  wire                uSystolicPE_423_io_clear_w_d;
  wire                uSystolicPE_423_io_enable_o_d;
  wire                uSystolicPE_423_io_clear_o_d;
  wire                uSystolicPE_423_io_ifm_sign_d;
  wire                uSystolicPE_423_io_ifm_dff_d;
  wire                uSystolicPE_423_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_423_io_randW_d;
  wire       [14:0]   uSystolicPE_423_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_423_io_ofm_d;
  wire                uSystolicPE_424_io_mac_done_d;
  wire                uSystolicPE_424_io_enable_i_d;
  wire                uSystolicPE_424_io_clear_i_d;
  wire                uSystolicPE_424_io_enable_w_d;
  wire                uSystolicPE_424_io_clear_w_d;
  wire                uSystolicPE_424_io_enable_o_d;
  wire                uSystolicPE_424_io_clear_o_d;
  wire                uSystolicPE_424_io_ifm_sign_d;
  wire                uSystolicPE_424_io_ifm_dff_d;
  wire                uSystolicPE_424_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_424_io_randW_d;
  wire       [14:0]   uSystolicPE_424_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_424_io_ofm_d;
  wire                uSystolicPE_425_io_mac_done_d;
  wire                uSystolicPE_425_io_enable_i_d;
  wire                uSystolicPE_425_io_clear_i_d;
  wire                uSystolicPE_425_io_enable_w_d;
  wire                uSystolicPE_425_io_clear_w_d;
  wire                uSystolicPE_425_io_enable_o_d;
  wire                uSystolicPE_425_io_clear_o_d;
  wire                uSystolicPE_425_io_ifm_sign_d;
  wire                uSystolicPE_425_io_ifm_dff_d;
  wire                uSystolicPE_425_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_425_io_randW_d;
  wire       [14:0]   uSystolicPE_425_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_425_io_ofm_d;
  wire                uSystolicPE_426_io_mac_done_d;
  wire                uSystolicPE_426_io_enable_i_d;
  wire                uSystolicPE_426_io_clear_i_d;
  wire                uSystolicPE_426_io_enable_w_d;
  wire                uSystolicPE_426_io_clear_w_d;
  wire                uSystolicPE_426_io_enable_o_d;
  wire                uSystolicPE_426_io_clear_o_d;
  wire                uSystolicPE_426_io_ifm_sign_d;
  wire                uSystolicPE_426_io_ifm_dff_d;
  wire                uSystolicPE_426_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_426_io_randW_d;
  wire       [14:0]   uSystolicPE_426_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_426_io_ofm_d;
  wire                uSystolicPE_427_io_mac_done_d;
  wire                uSystolicPE_427_io_enable_i_d;
  wire                uSystolicPE_427_io_clear_i_d;
  wire                uSystolicPE_427_io_enable_w_d;
  wire                uSystolicPE_427_io_clear_w_d;
  wire                uSystolicPE_427_io_enable_o_d;
  wire                uSystolicPE_427_io_clear_o_d;
  wire                uSystolicPE_427_io_ifm_sign_d;
  wire                uSystolicPE_427_io_ifm_dff_d;
  wire                uSystolicPE_427_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_427_io_randW_d;
  wire       [14:0]   uSystolicPE_427_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_427_io_ofm_d;
  wire                uSystolicPE_428_io_mac_done_d;
  wire                uSystolicPE_428_io_enable_i_d;
  wire                uSystolicPE_428_io_clear_i_d;
  wire                uSystolicPE_428_io_enable_w_d;
  wire                uSystolicPE_428_io_clear_w_d;
  wire                uSystolicPE_428_io_enable_o_d;
  wire                uSystolicPE_428_io_clear_o_d;
  wire                uSystolicPE_428_io_ifm_sign_d;
  wire                uSystolicPE_428_io_ifm_dff_d;
  wire                uSystolicPE_428_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_428_io_randW_d;
  wire       [14:0]   uSystolicPE_428_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_428_io_ofm_d;
  wire                uSystolicPE_429_io_mac_done_d;
  wire                uSystolicPE_429_io_enable_i_d;
  wire                uSystolicPE_429_io_clear_i_d;
  wire                uSystolicPE_429_io_enable_w_d;
  wire                uSystolicPE_429_io_clear_w_d;
  wire                uSystolicPE_429_io_enable_o_d;
  wire                uSystolicPE_429_io_clear_o_d;
  wire                uSystolicPE_429_io_ifm_sign_d;
  wire                uSystolicPE_429_io_ifm_dff_d;
  wire                uSystolicPE_429_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_429_io_randW_d;
  wire       [14:0]   uSystolicPE_429_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_429_io_ofm_d;
  wire                uSystolicPE_430_io_mac_done_d;
  wire                uSystolicPE_430_io_enable_i_d;
  wire                uSystolicPE_430_io_clear_i_d;
  wire                uSystolicPE_430_io_enable_w_d;
  wire                uSystolicPE_430_io_clear_w_d;
  wire                uSystolicPE_430_io_enable_o_d;
  wire                uSystolicPE_430_io_clear_o_d;
  wire                uSystolicPE_430_io_ifm_sign_d;
  wire                uSystolicPE_430_io_ifm_dff_d;
  wire                uSystolicPE_430_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_430_io_randW_d;
  wire       [14:0]   uSystolicPE_430_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_430_io_ofm_d;
  wire                uSystolicPE_431_io_mac_done_d;
  wire                uSystolicPE_431_io_enable_i_d;
  wire                uSystolicPE_431_io_clear_i_d;
  wire                uSystolicPE_431_io_enable_w_d;
  wire                uSystolicPE_431_io_clear_w_d;
  wire                uSystolicPE_431_io_enable_o_d;
  wire                uSystolicPE_431_io_clear_o_d;
  wire                uSystolicPE_431_io_ifm_sign_d;
  wire                uSystolicPE_431_io_ifm_dff_d;
  wire                uSystolicPE_431_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_431_io_randW_d;
  wire       [14:0]   uSystolicPE_431_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_431_io_ofm_d;
  wire                uSystolicPE_432_io_mac_done_d;
  wire                uSystolicPE_432_io_enable_i_d;
  wire                uSystolicPE_432_io_clear_i_d;
  wire                uSystolicPE_432_io_enable_w_d;
  wire                uSystolicPE_432_io_clear_w_d;
  wire                uSystolicPE_432_io_enable_o_d;
  wire                uSystolicPE_432_io_clear_o_d;
  wire                uSystolicPE_432_io_ifm_sign_d;
  wire                uSystolicPE_432_io_ifm_dff_d;
  wire                uSystolicPE_432_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_432_io_randW_d;
  wire       [14:0]   uSystolicPE_432_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_432_io_ofm_d;
  wire                uSystolicPE_433_io_mac_done_d;
  wire                uSystolicPE_433_io_enable_i_d;
  wire                uSystolicPE_433_io_clear_i_d;
  wire                uSystolicPE_433_io_enable_w_d;
  wire                uSystolicPE_433_io_clear_w_d;
  wire                uSystolicPE_433_io_enable_o_d;
  wire                uSystolicPE_433_io_clear_o_d;
  wire                uSystolicPE_433_io_ifm_sign_d;
  wire                uSystolicPE_433_io_ifm_dff_d;
  wire                uSystolicPE_433_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_433_io_randW_d;
  wire       [14:0]   uSystolicPE_433_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_433_io_ofm_d;
  wire                uSystolicPE_434_io_mac_done_d;
  wire                uSystolicPE_434_io_enable_i_d;
  wire                uSystolicPE_434_io_clear_i_d;
  wire                uSystolicPE_434_io_enable_w_d;
  wire                uSystolicPE_434_io_clear_w_d;
  wire                uSystolicPE_434_io_enable_o_d;
  wire                uSystolicPE_434_io_clear_o_d;
  wire                uSystolicPE_434_io_ifm_sign_d;
  wire                uSystolicPE_434_io_ifm_dff_d;
  wire                uSystolicPE_434_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_434_io_randW_d;
  wire       [14:0]   uSystolicPE_434_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_434_io_ofm_d;
  wire                uSystolicPEBorder_29_io_mac_done_d;
  wire                uSystolicPEBorder_29_io_enable_i_d;
  wire                uSystolicPEBorder_29_io_clear_i_d;
  wire                uSystolicPEBorder_29_io_enable_w_d;
  wire                uSystolicPEBorder_29_io_clear_w_d;
  wire                uSystolicPEBorder_29_io_enable_o_d;
  wire                uSystolicPEBorder_29_io_clear_o_d;
  wire                uSystolicPEBorder_29_io_ifm_sign_d;
  wire                uSystolicPEBorder_29_io_ifm_dff_d;
  wire                uSystolicPEBorder_29_io_wght_sign_d;
  wire       [14:0]   uSystolicPEBorder_29_io_randW_d;
  wire       [14:0]   uSystolicPEBorder_29_io_wght_abs_d;
  wire       [31:0]   uSystolicPEBorder_29_io_ofm_d;
  wire                uSystolicPE_435_io_mac_done_d;
  wire                uSystolicPE_435_io_enable_i_d;
  wire                uSystolicPE_435_io_clear_i_d;
  wire                uSystolicPE_435_io_enable_w_d;
  wire                uSystolicPE_435_io_clear_w_d;
  wire                uSystolicPE_435_io_enable_o_d;
  wire                uSystolicPE_435_io_clear_o_d;
  wire                uSystolicPE_435_io_ifm_sign_d;
  wire                uSystolicPE_435_io_ifm_dff_d;
  wire                uSystolicPE_435_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_435_io_randW_d;
  wire       [14:0]   uSystolicPE_435_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_435_io_ofm_d;
  wire                uSystolicPE_436_io_mac_done_d;
  wire                uSystolicPE_436_io_enable_i_d;
  wire                uSystolicPE_436_io_clear_i_d;
  wire                uSystolicPE_436_io_enable_w_d;
  wire                uSystolicPE_436_io_clear_w_d;
  wire                uSystolicPE_436_io_enable_o_d;
  wire                uSystolicPE_436_io_clear_o_d;
  wire                uSystolicPE_436_io_ifm_sign_d;
  wire                uSystolicPE_436_io_ifm_dff_d;
  wire                uSystolicPE_436_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_436_io_randW_d;
  wire       [14:0]   uSystolicPE_436_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_436_io_ofm_d;
  wire                uSystolicPE_437_io_mac_done_d;
  wire                uSystolicPE_437_io_enable_i_d;
  wire                uSystolicPE_437_io_clear_i_d;
  wire                uSystolicPE_437_io_enable_w_d;
  wire                uSystolicPE_437_io_clear_w_d;
  wire                uSystolicPE_437_io_enable_o_d;
  wire                uSystolicPE_437_io_clear_o_d;
  wire                uSystolicPE_437_io_ifm_sign_d;
  wire                uSystolicPE_437_io_ifm_dff_d;
  wire                uSystolicPE_437_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_437_io_randW_d;
  wire       [14:0]   uSystolicPE_437_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_437_io_ofm_d;
  wire                uSystolicPE_438_io_mac_done_d;
  wire                uSystolicPE_438_io_enable_i_d;
  wire                uSystolicPE_438_io_clear_i_d;
  wire                uSystolicPE_438_io_enable_w_d;
  wire                uSystolicPE_438_io_clear_w_d;
  wire                uSystolicPE_438_io_enable_o_d;
  wire                uSystolicPE_438_io_clear_o_d;
  wire                uSystolicPE_438_io_ifm_sign_d;
  wire                uSystolicPE_438_io_ifm_dff_d;
  wire                uSystolicPE_438_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_438_io_randW_d;
  wire       [14:0]   uSystolicPE_438_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_438_io_ofm_d;
  wire                uSystolicPE_439_io_mac_done_d;
  wire                uSystolicPE_439_io_enable_i_d;
  wire                uSystolicPE_439_io_clear_i_d;
  wire                uSystolicPE_439_io_enable_w_d;
  wire                uSystolicPE_439_io_clear_w_d;
  wire                uSystolicPE_439_io_enable_o_d;
  wire                uSystolicPE_439_io_clear_o_d;
  wire                uSystolicPE_439_io_ifm_sign_d;
  wire                uSystolicPE_439_io_ifm_dff_d;
  wire                uSystolicPE_439_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_439_io_randW_d;
  wire       [14:0]   uSystolicPE_439_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_439_io_ofm_d;
  wire                uSystolicPE_440_io_mac_done_d;
  wire                uSystolicPE_440_io_enable_i_d;
  wire                uSystolicPE_440_io_clear_i_d;
  wire                uSystolicPE_440_io_enable_w_d;
  wire                uSystolicPE_440_io_clear_w_d;
  wire                uSystolicPE_440_io_enable_o_d;
  wire                uSystolicPE_440_io_clear_o_d;
  wire                uSystolicPE_440_io_ifm_sign_d;
  wire                uSystolicPE_440_io_ifm_dff_d;
  wire                uSystolicPE_440_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_440_io_randW_d;
  wire       [14:0]   uSystolicPE_440_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_440_io_ofm_d;
  wire                uSystolicPE_441_io_mac_done_d;
  wire                uSystolicPE_441_io_enable_i_d;
  wire                uSystolicPE_441_io_clear_i_d;
  wire                uSystolicPE_441_io_enable_w_d;
  wire                uSystolicPE_441_io_clear_w_d;
  wire                uSystolicPE_441_io_enable_o_d;
  wire                uSystolicPE_441_io_clear_o_d;
  wire                uSystolicPE_441_io_ifm_sign_d;
  wire                uSystolicPE_441_io_ifm_dff_d;
  wire                uSystolicPE_441_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_441_io_randW_d;
  wire       [14:0]   uSystolicPE_441_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_441_io_ofm_d;
  wire                uSystolicPE_442_io_mac_done_d;
  wire                uSystolicPE_442_io_enable_i_d;
  wire                uSystolicPE_442_io_clear_i_d;
  wire                uSystolicPE_442_io_enable_w_d;
  wire                uSystolicPE_442_io_clear_w_d;
  wire                uSystolicPE_442_io_enable_o_d;
  wire                uSystolicPE_442_io_clear_o_d;
  wire                uSystolicPE_442_io_ifm_sign_d;
  wire                uSystolicPE_442_io_ifm_dff_d;
  wire                uSystolicPE_442_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_442_io_randW_d;
  wire       [14:0]   uSystolicPE_442_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_442_io_ofm_d;
  wire                uSystolicPE_443_io_mac_done_d;
  wire                uSystolicPE_443_io_enable_i_d;
  wire                uSystolicPE_443_io_clear_i_d;
  wire                uSystolicPE_443_io_enable_w_d;
  wire                uSystolicPE_443_io_clear_w_d;
  wire                uSystolicPE_443_io_enable_o_d;
  wire                uSystolicPE_443_io_clear_o_d;
  wire                uSystolicPE_443_io_ifm_sign_d;
  wire                uSystolicPE_443_io_ifm_dff_d;
  wire                uSystolicPE_443_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_443_io_randW_d;
  wire       [14:0]   uSystolicPE_443_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_443_io_ofm_d;
  wire                uSystolicPE_444_io_mac_done_d;
  wire                uSystolicPE_444_io_enable_i_d;
  wire                uSystolicPE_444_io_clear_i_d;
  wire                uSystolicPE_444_io_enable_w_d;
  wire                uSystolicPE_444_io_clear_w_d;
  wire                uSystolicPE_444_io_enable_o_d;
  wire                uSystolicPE_444_io_clear_o_d;
  wire                uSystolicPE_444_io_ifm_sign_d;
  wire                uSystolicPE_444_io_ifm_dff_d;
  wire                uSystolicPE_444_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_444_io_randW_d;
  wire       [14:0]   uSystolicPE_444_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_444_io_ofm_d;
  wire                uSystolicPE_445_io_mac_done_d;
  wire                uSystolicPE_445_io_enable_i_d;
  wire                uSystolicPE_445_io_clear_i_d;
  wire                uSystolicPE_445_io_enable_w_d;
  wire                uSystolicPE_445_io_clear_w_d;
  wire                uSystolicPE_445_io_enable_o_d;
  wire                uSystolicPE_445_io_clear_o_d;
  wire                uSystolicPE_445_io_ifm_sign_d;
  wire                uSystolicPE_445_io_ifm_dff_d;
  wire                uSystolicPE_445_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_445_io_randW_d;
  wire       [14:0]   uSystolicPE_445_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_445_io_ofm_d;
  wire                uSystolicPE_446_io_mac_done_d;
  wire                uSystolicPE_446_io_enable_i_d;
  wire                uSystolicPE_446_io_clear_i_d;
  wire                uSystolicPE_446_io_enable_w_d;
  wire                uSystolicPE_446_io_clear_w_d;
  wire                uSystolicPE_446_io_enable_o_d;
  wire                uSystolicPE_446_io_clear_o_d;
  wire                uSystolicPE_446_io_ifm_sign_d;
  wire                uSystolicPE_446_io_ifm_dff_d;
  wire                uSystolicPE_446_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_446_io_randW_d;
  wire       [14:0]   uSystolicPE_446_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_446_io_ofm_d;
  wire                uSystolicPE_447_io_mac_done_d;
  wire                uSystolicPE_447_io_enable_i_d;
  wire                uSystolicPE_447_io_clear_i_d;
  wire                uSystolicPE_447_io_enable_w_d;
  wire                uSystolicPE_447_io_clear_w_d;
  wire                uSystolicPE_447_io_enable_o_d;
  wire                uSystolicPE_447_io_clear_o_d;
  wire                uSystolicPE_447_io_ifm_sign_d;
  wire                uSystolicPE_447_io_ifm_dff_d;
  wire                uSystolicPE_447_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_447_io_randW_d;
  wire       [14:0]   uSystolicPE_447_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_447_io_ofm_d;
  wire                uSystolicPE_448_io_mac_done_d;
  wire                uSystolicPE_448_io_enable_i_d;
  wire                uSystolicPE_448_io_clear_i_d;
  wire                uSystolicPE_448_io_enable_w_d;
  wire                uSystolicPE_448_io_clear_w_d;
  wire                uSystolicPE_448_io_enable_o_d;
  wire                uSystolicPE_448_io_clear_o_d;
  wire                uSystolicPE_448_io_ifm_sign_d;
  wire                uSystolicPE_448_io_ifm_dff_d;
  wire                uSystolicPE_448_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_448_io_randW_d;
  wire       [14:0]   uSystolicPE_448_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_448_io_ofm_d;
  wire                uSystolicPE_449_io_mac_done_d;
  wire                uSystolicPE_449_io_enable_i_d;
  wire                uSystolicPE_449_io_clear_i_d;
  wire                uSystolicPE_449_io_enable_w_d;
  wire                uSystolicPE_449_io_clear_w_d;
  wire                uSystolicPE_449_io_enable_o_d;
  wire                uSystolicPE_449_io_clear_o_d;
  wire                uSystolicPE_449_io_ifm_sign_d;
  wire                uSystolicPE_449_io_ifm_dff_d;
  wire                uSystolicPE_449_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_449_io_randW_d;
  wire       [14:0]   uSystolicPE_449_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_449_io_ofm_d;
  wire                uSystolicPEBorder_30_io_mac_done_d;
  wire                uSystolicPEBorder_30_io_enable_i_d;
  wire                uSystolicPEBorder_30_io_clear_i_d;
  wire                uSystolicPEBorder_30_io_enable_w_d;
  wire                uSystolicPEBorder_30_io_clear_w_d;
  wire                uSystolicPEBorder_30_io_enable_o_d;
  wire                uSystolicPEBorder_30_io_clear_o_d;
  wire                uSystolicPEBorder_30_io_ifm_sign_d;
  wire                uSystolicPEBorder_30_io_ifm_dff_d;
  wire                uSystolicPEBorder_30_io_wght_sign_d;
  wire       [14:0]   uSystolicPEBorder_30_io_randW_d;
  wire       [14:0]   uSystolicPEBorder_30_io_wght_abs_d;
  wire       [31:0]   uSystolicPEBorder_30_io_ofm_d;
  wire                uSystolicPE_450_io_mac_done_d;
  wire                uSystolicPE_450_io_enable_i_d;
  wire                uSystolicPE_450_io_clear_i_d;
  wire                uSystolicPE_450_io_enable_w_d;
  wire                uSystolicPE_450_io_clear_w_d;
  wire                uSystolicPE_450_io_enable_o_d;
  wire                uSystolicPE_450_io_clear_o_d;
  wire                uSystolicPE_450_io_ifm_sign_d;
  wire                uSystolicPE_450_io_ifm_dff_d;
  wire                uSystolicPE_450_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_450_io_randW_d;
  wire       [14:0]   uSystolicPE_450_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_450_io_ofm_d;
  wire                uSystolicPE_451_io_mac_done_d;
  wire                uSystolicPE_451_io_enable_i_d;
  wire                uSystolicPE_451_io_clear_i_d;
  wire                uSystolicPE_451_io_enable_w_d;
  wire                uSystolicPE_451_io_clear_w_d;
  wire                uSystolicPE_451_io_enable_o_d;
  wire                uSystolicPE_451_io_clear_o_d;
  wire                uSystolicPE_451_io_ifm_sign_d;
  wire                uSystolicPE_451_io_ifm_dff_d;
  wire                uSystolicPE_451_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_451_io_randW_d;
  wire       [14:0]   uSystolicPE_451_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_451_io_ofm_d;
  wire                uSystolicPE_452_io_mac_done_d;
  wire                uSystolicPE_452_io_enable_i_d;
  wire                uSystolicPE_452_io_clear_i_d;
  wire                uSystolicPE_452_io_enable_w_d;
  wire                uSystolicPE_452_io_clear_w_d;
  wire                uSystolicPE_452_io_enable_o_d;
  wire                uSystolicPE_452_io_clear_o_d;
  wire                uSystolicPE_452_io_ifm_sign_d;
  wire                uSystolicPE_452_io_ifm_dff_d;
  wire                uSystolicPE_452_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_452_io_randW_d;
  wire       [14:0]   uSystolicPE_452_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_452_io_ofm_d;
  wire                uSystolicPE_453_io_mac_done_d;
  wire                uSystolicPE_453_io_enable_i_d;
  wire                uSystolicPE_453_io_clear_i_d;
  wire                uSystolicPE_453_io_enable_w_d;
  wire                uSystolicPE_453_io_clear_w_d;
  wire                uSystolicPE_453_io_enable_o_d;
  wire                uSystolicPE_453_io_clear_o_d;
  wire                uSystolicPE_453_io_ifm_sign_d;
  wire                uSystolicPE_453_io_ifm_dff_d;
  wire                uSystolicPE_453_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_453_io_randW_d;
  wire       [14:0]   uSystolicPE_453_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_453_io_ofm_d;
  wire                uSystolicPE_454_io_mac_done_d;
  wire                uSystolicPE_454_io_enable_i_d;
  wire                uSystolicPE_454_io_clear_i_d;
  wire                uSystolicPE_454_io_enable_w_d;
  wire                uSystolicPE_454_io_clear_w_d;
  wire                uSystolicPE_454_io_enable_o_d;
  wire                uSystolicPE_454_io_clear_o_d;
  wire                uSystolicPE_454_io_ifm_sign_d;
  wire                uSystolicPE_454_io_ifm_dff_d;
  wire                uSystolicPE_454_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_454_io_randW_d;
  wire       [14:0]   uSystolicPE_454_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_454_io_ofm_d;
  wire                uSystolicPE_455_io_mac_done_d;
  wire                uSystolicPE_455_io_enable_i_d;
  wire                uSystolicPE_455_io_clear_i_d;
  wire                uSystolicPE_455_io_enable_w_d;
  wire                uSystolicPE_455_io_clear_w_d;
  wire                uSystolicPE_455_io_enable_o_d;
  wire                uSystolicPE_455_io_clear_o_d;
  wire                uSystolicPE_455_io_ifm_sign_d;
  wire                uSystolicPE_455_io_ifm_dff_d;
  wire                uSystolicPE_455_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_455_io_randW_d;
  wire       [14:0]   uSystolicPE_455_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_455_io_ofm_d;
  wire                uSystolicPE_456_io_mac_done_d;
  wire                uSystolicPE_456_io_enable_i_d;
  wire                uSystolicPE_456_io_clear_i_d;
  wire                uSystolicPE_456_io_enable_w_d;
  wire                uSystolicPE_456_io_clear_w_d;
  wire                uSystolicPE_456_io_enable_o_d;
  wire                uSystolicPE_456_io_clear_o_d;
  wire                uSystolicPE_456_io_ifm_sign_d;
  wire                uSystolicPE_456_io_ifm_dff_d;
  wire                uSystolicPE_456_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_456_io_randW_d;
  wire       [14:0]   uSystolicPE_456_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_456_io_ofm_d;
  wire                uSystolicPE_457_io_mac_done_d;
  wire                uSystolicPE_457_io_enable_i_d;
  wire                uSystolicPE_457_io_clear_i_d;
  wire                uSystolicPE_457_io_enable_w_d;
  wire                uSystolicPE_457_io_clear_w_d;
  wire                uSystolicPE_457_io_enable_o_d;
  wire                uSystolicPE_457_io_clear_o_d;
  wire                uSystolicPE_457_io_ifm_sign_d;
  wire                uSystolicPE_457_io_ifm_dff_d;
  wire                uSystolicPE_457_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_457_io_randW_d;
  wire       [14:0]   uSystolicPE_457_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_457_io_ofm_d;
  wire                uSystolicPE_458_io_mac_done_d;
  wire                uSystolicPE_458_io_enable_i_d;
  wire                uSystolicPE_458_io_clear_i_d;
  wire                uSystolicPE_458_io_enable_w_d;
  wire                uSystolicPE_458_io_clear_w_d;
  wire                uSystolicPE_458_io_enable_o_d;
  wire                uSystolicPE_458_io_clear_o_d;
  wire                uSystolicPE_458_io_ifm_sign_d;
  wire                uSystolicPE_458_io_ifm_dff_d;
  wire                uSystolicPE_458_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_458_io_randW_d;
  wire       [14:0]   uSystolicPE_458_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_458_io_ofm_d;
  wire                uSystolicPE_459_io_mac_done_d;
  wire                uSystolicPE_459_io_enable_i_d;
  wire                uSystolicPE_459_io_clear_i_d;
  wire                uSystolicPE_459_io_enable_w_d;
  wire                uSystolicPE_459_io_clear_w_d;
  wire                uSystolicPE_459_io_enable_o_d;
  wire                uSystolicPE_459_io_clear_o_d;
  wire                uSystolicPE_459_io_ifm_sign_d;
  wire                uSystolicPE_459_io_ifm_dff_d;
  wire                uSystolicPE_459_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_459_io_randW_d;
  wire       [14:0]   uSystolicPE_459_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_459_io_ofm_d;
  wire                uSystolicPE_460_io_mac_done_d;
  wire                uSystolicPE_460_io_enable_i_d;
  wire                uSystolicPE_460_io_clear_i_d;
  wire                uSystolicPE_460_io_enable_w_d;
  wire                uSystolicPE_460_io_clear_w_d;
  wire                uSystolicPE_460_io_enable_o_d;
  wire                uSystolicPE_460_io_clear_o_d;
  wire                uSystolicPE_460_io_ifm_sign_d;
  wire                uSystolicPE_460_io_ifm_dff_d;
  wire                uSystolicPE_460_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_460_io_randW_d;
  wire       [14:0]   uSystolicPE_460_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_460_io_ofm_d;
  wire                uSystolicPE_461_io_mac_done_d;
  wire                uSystolicPE_461_io_enable_i_d;
  wire                uSystolicPE_461_io_clear_i_d;
  wire                uSystolicPE_461_io_enable_w_d;
  wire                uSystolicPE_461_io_clear_w_d;
  wire                uSystolicPE_461_io_enable_o_d;
  wire                uSystolicPE_461_io_clear_o_d;
  wire                uSystolicPE_461_io_ifm_sign_d;
  wire                uSystolicPE_461_io_ifm_dff_d;
  wire                uSystolicPE_461_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_461_io_randW_d;
  wire       [14:0]   uSystolicPE_461_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_461_io_ofm_d;
  wire                uSystolicPE_462_io_mac_done_d;
  wire                uSystolicPE_462_io_enable_i_d;
  wire                uSystolicPE_462_io_clear_i_d;
  wire                uSystolicPE_462_io_enable_w_d;
  wire                uSystolicPE_462_io_clear_w_d;
  wire                uSystolicPE_462_io_enable_o_d;
  wire                uSystolicPE_462_io_clear_o_d;
  wire                uSystolicPE_462_io_ifm_sign_d;
  wire                uSystolicPE_462_io_ifm_dff_d;
  wire                uSystolicPE_462_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_462_io_randW_d;
  wire       [14:0]   uSystolicPE_462_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_462_io_ofm_d;
  wire                uSystolicPE_463_io_mac_done_d;
  wire                uSystolicPE_463_io_enable_i_d;
  wire                uSystolicPE_463_io_clear_i_d;
  wire                uSystolicPE_463_io_enable_w_d;
  wire                uSystolicPE_463_io_clear_w_d;
  wire                uSystolicPE_463_io_enable_o_d;
  wire                uSystolicPE_463_io_clear_o_d;
  wire                uSystolicPE_463_io_ifm_sign_d;
  wire                uSystolicPE_463_io_ifm_dff_d;
  wire                uSystolicPE_463_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_463_io_randW_d;
  wire       [14:0]   uSystolicPE_463_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_463_io_ofm_d;
  wire                uSystolicPE_464_io_mac_done_d;
  wire                uSystolicPE_464_io_enable_i_d;
  wire                uSystolicPE_464_io_clear_i_d;
  wire                uSystolicPE_464_io_enable_w_d;
  wire                uSystolicPE_464_io_clear_w_d;
  wire                uSystolicPE_464_io_enable_o_d;
  wire                uSystolicPE_464_io_clear_o_d;
  wire                uSystolicPE_464_io_ifm_sign_d;
  wire                uSystolicPE_464_io_ifm_dff_d;
  wire                uSystolicPE_464_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_464_io_randW_d;
  wire       [14:0]   uSystolicPE_464_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_464_io_ofm_d;
  wire                uSystolicPEBorder_31_io_mac_done_d;
  wire                uSystolicPEBorder_31_io_enable_i_d;
  wire                uSystolicPEBorder_31_io_clear_i_d;
  wire                uSystolicPEBorder_31_io_enable_w_d;
  wire                uSystolicPEBorder_31_io_clear_w_d;
  wire                uSystolicPEBorder_31_io_enable_o_d;
  wire                uSystolicPEBorder_31_io_clear_o_d;
  wire                uSystolicPEBorder_31_io_ifm_sign_d;
  wire                uSystolicPEBorder_31_io_ifm_dff_d;
  wire                uSystolicPEBorder_31_io_wght_sign_d;
  wire       [14:0]   uSystolicPEBorder_31_io_randW_d;
  wire       [14:0]   uSystolicPEBorder_31_io_wght_abs_d;
  wire       [31:0]   uSystolicPEBorder_31_io_ofm_d;
  wire                uSystolicPE_465_io_mac_done_d;
  wire                uSystolicPE_465_io_enable_i_d;
  wire                uSystolicPE_465_io_clear_i_d;
  wire                uSystolicPE_465_io_enable_w_d;
  wire                uSystolicPE_465_io_clear_w_d;
  wire                uSystolicPE_465_io_enable_o_d;
  wire                uSystolicPE_465_io_clear_o_d;
  wire                uSystolicPE_465_io_ifm_sign_d;
  wire                uSystolicPE_465_io_ifm_dff_d;
  wire                uSystolicPE_465_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_465_io_randW_d;
  wire       [14:0]   uSystolicPE_465_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_465_io_ofm_d;
  wire                uSystolicPE_466_io_mac_done_d;
  wire                uSystolicPE_466_io_enable_i_d;
  wire                uSystolicPE_466_io_clear_i_d;
  wire                uSystolicPE_466_io_enable_w_d;
  wire                uSystolicPE_466_io_clear_w_d;
  wire                uSystolicPE_466_io_enable_o_d;
  wire                uSystolicPE_466_io_clear_o_d;
  wire                uSystolicPE_466_io_ifm_sign_d;
  wire                uSystolicPE_466_io_ifm_dff_d;
  wire                uSystolicPE_466_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_466_io_randW_d;
  wire       [14:0]   uSystolicPE_466_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_466_io_ofm_d;
  wire                uSystolicPE_467_io_mac_done_d;
  wire                uSystolicPE_467_io_enable_i_d;
  wire                uSystolicPE_467_io_clear_i_d;
  wire                uSystolicPE_467_io_enable_w_d;
  wire                uSystolicPE_467_io_clear_w_d;
  wire                uSystolicPE_467_io_enable_o_d;
  wire                uSystolicPE_467_io_clear_o_d;
  wire                uSystolicPE_467_io_ifm_sign_d;
  wire                uSystolicPE_467_io_ifm_dff_d;
  wire                uSystolicPE_467_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_467_io_randW_d;
  wire       [14:0]   uSystolicPE_467_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_467_io_ofm_d;
  wire                uSystolicPE_468_io_mac_done_d;
  wire                uSystolicPE_468_io_enable_i_d;
  wire                uSystolicPE_468_io_clear_i_d;
  wire                uSystolicPE_468_io_enable_w_d;
  wire                uSystolicPE_468_io_clear_w_d;
  wire                uSystolicPE_468_io_enable_o_d;
  wire                uSystolicPE_468_io_clear_o_d;
  wire                uSystolicPE_468_io_ifm_sign_d;
  wire                uSystolicPE_468_io_ifm_dff_d;
  wire                uSystolicPE_468_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_468_io_randW_d;
  wire       [14:0]   uSystolicPE_468_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_468_io_ofm_d;
  wire                uSystolicPE_469_io_mac_done_d;
  wire                uSystolicPE_469_io_enable_i_d;
  wire                uSystolicPE_469_io_clear_i_d;
  wire                uSystolicPE_469_io_enable_w_d;
  wire                uSystolicPE_469_io_clear_w_d;
  wire                uSystolicPE_469_io_enable_o_d;
  wire                uSystolicPE_469_io_clear_o_d;
  wire                uSystolicPE_469_io_ifm_sign_d;
  wire                uSystolicPE_469_io_ifm_dff_d;
  wire                uSystolicPE_469_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_469_io_randW_d;
  wire       [14:0]   uSystolicPE_469_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_469_io_ofm_d;
  wire                uSystolicPE_470_io_mac_done_d;
  wire                uSystolicPE_470_io_enable_i_d;
  wire                uSystolicPE_470_io_clear_i_d;
  wire                uSystolicPE_470_io_enable_w_d;
  wire                uSystolicPE_470_io_clear_w_d;
  wire                uSystolicPE_470_io_enable_o_d;
  wire                uSystolicPE_470_io_clear_o_d;
  wire                uSystolicPE_470_io_ifm_sign_d;
  wire                uSystolicPE_470_io_ifm_dff_d;
  wire                uSystolicPE_470_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_470_io_randW_d;
  wire       [14:0]   uSystolicPE_470_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_470_io_ofm_d;
  wire                uSystolicPE_471_io_mac_done_d;
  wire                uSystolicPE_471_io_enable_i_d;
  wire                uSystolicPE_471_io_clear_i_d;
  wire                uSystolicPE_471_io_enable_w_d;
  wire                uSystolicPE_471_io_clear_w_d;
  wire                uSystolicPE_471_io_enable_o_d;
  wire                uSystolicPE_471_io_clear_o_d;
  wire                uSystolicPE_471_io_ifm_sign_d;
  wire                uSystolicPE_471_io_ifm_dff_d;
  wire                uSystolicPE_471_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_471_io_randW_d;
  wire       [14:0]   uSystolicPE_471_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_471_io_ofm_d;
  wire                uSystolicPE_472_io_mac_done_d;
  wire                uSystolicPE_472_io_enable_i_d;
  wire                uSystolicPE_472_io_clear_i_d;
  wire                uSystolicPE_472_io_enable_w_d;
  wire                uSystolicPE_472_io_clear_w_d;
  wire                uSystolicPE_472_io_enable_o_d;
  wire                uSystolicPE_472_io_clear_o_d;
  wire                uSystolicPE_472_io_ifm_sign_d;
  wire                uSystolicPE_472_io_ifm_dff_d;
  wire                uSystolicPE_472_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_472_io_randW_d;
  wire       [14:0]   uSystolicPE_472_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_472_io_ofm_d;
  wire                uSystolicPE_473_io_mac_done_d;
  wire                uSystolicPE_473_io_enable_i_d;
  wire                uSystolicPE_473_io_clear_i_d;
  wire                uSystolicPE_473_io_enable_w_d;
  wire                uSystolicPE_473_io_clear_w_d;
  wire                uSystolicPE_473_io_enable_o_d;
  wire                uSystolicPE_473_io_clear_o_d;
  wire                uSystolicPE_473_io_ifm_sign_d;
  wire                uSystolicPE_473_io_ifm_dff_d;
  wire                uSystolicPE_473_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_473_io_randW_d;
  wire       [14:0]   uSystolicPE_473_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_473_io_ofm_d;
  wire                uSystolicPE_474_io_mac_done_d;
  wire                uSystolicPE_474_io_enable_i_d;
  wire                uSystolicPE_474_io_clear_i_d;
  wire                uSystolicPE_474_io_enable_w_d;
  wire                uSystolicPE_474_io_clear_w_d;
  wire                uSystolicPE_474_io_enable_o_d;
  wire                uSystolicPE_474_io_clear_o_d;
  wire                uSystolicPE_474_io_ifm_sign_d;
  wire                uSystolicPE_474_io_ifm_dff_d;
  wire                uSystolicPE_474_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_474_io_randW_d;
  wire       [14:0]   uSystolicPE_474_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_474_io_ofm_d;
  wire                uSystolicPE_475_io_mac_done_d;
  wire                uSystolicPE_475_io_enable_i_d;
  wire                uSystolicPE_475_io_clear_i_d;
  wire                uSystolicPE_475_io_enable_w_d;
  wire                uSystolicPE_475_io_clear_w_d;
  wire                uSystolicPE_475_io_enable_o_d;
  wire                uSystolicPE_475_io_clear_o_d;
  wire                uSystolicPE_475_io_ifm_sign_d;
  wire                uSystolicPE_475_io_ifm_dff_d;
  wire                uSystolicPE_475_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_475_io_randW_d;
  wire       [14:0]   uSystolicPE_475_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_475_io_ofm_d;
  wire                uSystolicPE_476_io_mac_done_d;
  wire                uSystolicPE_476_io_enable_i_d;
  wire                uSystolicPE_476_io_clear_i_d;
  wire                uSystolicPE_476_io_enable_w_d;
  wire                uSystolicPE_476_io_clear_w_d;
  wire                uSystolicPE_476_io_enable_o_d;
  wire                uSystolicPE_476_io_clear_o_d;
  wire                uSystolicPE_476_io_ifm_sign_d;
  wire                uSystolicPE_476_io_ifm_dff_d;
  wire                uSystolicPE_476_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_476_io_randW_d;
  wire       [14:0]   uSystolicPE_476_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_476_io_ofm_d;
  wire                uSystolicPE_477_io_mac_done_d;
  wire                uSystolicPE_477_io_enable_i_d;
  wire                uSystolicPE_477_io_clear_i_d;
  wire                uSystolicPE_477_io_enable_w_d;
  wire                uSystolicPE_477_io_clear_w_d;
  wire                uSystolicPE_477_io_enable_o_d;
  wire                uSystolicPE_477_io_clear_o_d;
  wire                uSystolicPE_477_io_ifm_sign_d;
  wire                uSystolicPE_477_io_ifm_dff_d;
  wire                uSystolicPE_477_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_477_io_randW_d;
  wire       [14:0]   uSystolicPE_477_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_477_io_ofm_d;
  wire                uSystolicPE_478_io_mac_done_d;
  wire                uSystolicPE_478_io_enable_i_d;
  wire                uSystolicPE_478_io_clear_i_d;
  wire                uSystolicPE_478_io_enable_w_d;
  wire                uSystolicPE_478_io_clear_w_d;
  wire                uSystolicPE_478_io_enable_o_d;
  wire                uSystolicPE_478_io_clear_o_d;
  wire                uSystolicPE_478_io_ifm_sign_d;
  wire                uSystolicPE_478_io_ifm_dff_d;
  wire                uSystolicPE_478_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_478_io_randW_d;
  wire       [14:0]   uSystolicPE_478_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_478_io_ofm_d;
  wire                uSystolicPE_479_io_mac_done_d;
  wire                uSystolicPE_479_io_enable_i_d;
  wire                uSystolicPE_479_io_clear_i_d;
  wire                uSystolicPE_479_io_enable_w_d;
  wire                uSystolicPE_479_io_clear_w_d;
  wire                uSystolicPE_479_io_enable_o_d;
  wire                uSystolicPE_479_io_clear_o_d;
  wire                uSystolicPE_479_io_ifm_sign_d;
  wire                uSystolicPE_479_io_ifm_dff_d;
  wire                uSystolicPE_479_io_wght_sign_d;
  wire       [14:0]   uSystolicPE_479_io_randW_d;
  wire       [14:0]   uSystolicPE_479_io_wght_abs_d;
  wire       [31:0]   uSystolicPE_479_io_ofm_d;
  reg        [16:0]   enable_i_x_0;
  reg        [16:0]   enable_i_x_1;
  reg        [16:0]   enable_i_x_2;
  reg        [16:0]   enable_i_x_3;
  reg        [16:0]   enable_i_x_4;
  reg        [16:0]   enable_i_x_5;
  reg        [16:0]   enable_i_x_6;
  reg        [16:0]   enable_i_x_7;
  reg        [16:0]   enable_i_x_8;
  reg        [16:0]   enable_i_x_9;
  reg        [16:0]   enable_i_x_10;
  reg        [16:0]   enable_i_x_11;
  reg        [16:0]   enable_i_x_12;
  reg        [16:0]   enable_i_x_13;
  reg        [16:0]   enable_i_x_14;
  reg        [16:0]   enable_i_x_15;
  reg        [16:0]   clear_i_x_0;
  reg        [16:0]   clear_i_x_1;
  reg        [16:0]   clear_i_x_2;
  reg        [16:0]   clear_i_x_3;
  reg        [16:0]   clear_i_x_4;
  reg        [16:0]   clear_i_x_5;
  reg        [16:0]   clear_i_x_6;
  reg        [16:0]   clear_i_x_7;
  reg        [16:0]   clear_i_x_8;
  reg        [16:0]   clear_i_x_9;
  reg        [16:0]   clear_i_x_10;
  reg        [16:0]   clear_i_x_11;
  reg        [16:0]   clear_i_x_12;
  reg        [16:0]   clear_i_x_13;
  reg        [16:0]   clear_i_x_14;
  reg        [16:0]   clear_i_x_15;
  reg        [16:0]   mac_done_x_0;
  reg        [16:0]   mac_done_x_1;
  reg        [16:0]   mac_done_x_2;
  reg        [16:0]   mac_done_x_3;
  reg        [16:0]   mac_done_x_4;
  reg        [16:0]   mac_done_x_5;
  reg        [16:0]   mac_done_x_6;
  reg        [16:0]   mac_done_x_7;
  reg        [16:0]   mac_done_x_8;
  reg        [16:0]   mac_done_x_9;
  reg        [16:0]   mac_done_x_10;
  reg        [16:0]   mac_done_x_11;
  reg        [16:0]   mac_done_x_12;
  reg        [16:0]   mac_done_x_13;
  reg        [16:0]   mac_done_x_14;
  reg        [16:0]   mac_done_x_15;
  reg        [16:0]   enable_w_x_0;
  reg        [16:0]   enable_w_x_1;
  reg        [16:0]   enable_w_x_2;
  reg        [16:0]   enable_w_x_3;
  reg        [16:0]   enable_w_x_4;
  reg        [16:0]   enable_w_x_5;
  reg        [16:0]   enable_w_x_6;
  reg        [16:0]   enable_w_x_7;
  reg        [16:0]   enable_w_x_8;
  reg        [16:0]   enable_w_x_9;
  reg        [16:0]   enable_w_x_10;
  reg        [16:0]   enable_w_x_11;
  reg        [16:0]   enable_w_x_12;
  reg        [16:0]   enable_w_x_13;
  reg        [16:0]   enable_w_x_14;
  reg        [16:0]   enable_w_x_15;
  reg        [16:0]   clear_w_x_0;
  reg        [16:0]   clear_w_x_1;
  reg        [16:0]   clear_w_x_2;
  reg        [16:0]   clear_w_x_3;
  reg        [16:0]   clear_w_x_4;
  reg        [16:0]   clear_w_x_5;
  reg        [16:0]   clear_w_x_6;
  reg        [16:0]   clear_w_x_7;
  reg        [16:0]   clear_w_x_8;
  reg        [16:0]   clear_w_x_9;
  reg        [16:0]   clear_w_x_10;
  reg        [16:0]   clear_w_x_11;
  reg        [16:0]   clear_w_x_12;
  reg        [16:0]   clear_w_x_13;
  reg        [16:0]   clear_w_x_14;
  reg        [16:0]   clear_w_x_15;
  reg        [16:0]   enable_o_x_0;
  reg        [16:0]   enable_o_x_1;
  reg        [16:0]   enable_o_x_2;
  reg        [16:0]   enable_o_x_3;
  reg        [16:0]   enable_o_x_4;
  reg        [16:0]   enable_o_x_5;
  reg        [16:0]   enable_o_x_6;
  reg        [16:0]   enable_o_x_7;
  reg        [16:0]   enable_o_x_8;
  reg        [16:0]   enable_o_x_9;
  reg        [16:0]   enable_o_x_10;
  reg        [16:0]   enable_o_x_11;
  reg        [16:0]   enable_o_x_12;
  reg        [16:0]   enable_o_x_13;
  reg        [16:0]   enable_o_x_14;
  reg        [16:0]   enable_o_x_15;
  reg        [16:0]   clear_o_x_0;
  reg        [16:0]   clear_o_x_1;
  reg        [16:0]   clear_o_x_2;
  reg        [16:0]   clear_o_x_3;
  reg        [16:0]   clear_o_x_4;
  reg        [16:0]   clear_o_x_5;
  reg        [16:0]   clear_o_x_6;
  reg        [16:0]   clear_o_x_7;
  reg        [16:0]   clear_o_x_8;
  reg        [16:0]   clear_o_x_9;
  reg        [16:0]   clear_o_x_10;
  reg        [16:0]   clear_o_x_11;
  reg        [16:0]   clear_o_x_12;
  reg        [16:0]   clear_o_x_13;
  reg        [16:0]   clear_o_x_14;
  reg        [16:0]   clear_o_x_15;
  wire                ifm_sign_x_0_0;
  wire                ifm_sign_x_0_1;
  wire                ifm_sign_x_0_2;
  wire                ifm_sign_x_0_3;
  wire                ifm_sign_x_0_4;
  wire                ifm_sign_x_0_5;
  wire                ifm_sign_x_0_6;
  wire                ifm_sign_x_0_7;
  wire                ifm_sign_x_0_8;
  wire                ifm_sign_x_0_9;
  wire                ifm_sign_x_0_10;
  wire                ifm_sign_x_0_11;
  wire                ifm_sign_x_0_12;
  wire                ifm_sign_x_0_13;
  wire                ifm_sign_x_0_14;
  wire                ifm_sign_x_0_15;
  wire                ifm_sign_x_0_16;
  wire                ifm_sign_x_1_0;
  wire                ifm_sign_x_1_1;
  wire                ifm_sign_x_1_2;
  wire                ifm_sign_x_1_3;
  wire                ifm_sign_x_1_4;
  wire                ifm_sign_x_1_5;
  wire                ifm_sign_x_1_6;
  wire                ifm_sign_x_1_7;
  wire                ifm_sign_x_1_8;
  wire                ifm_sign_x_1_9;
  wire                ifm_sign_x_1_10;
  wire                ifm_sign_x_1_11;
  wire                ifm_sign_x_1_12;
  wire                ifm_sign_x_1_13;
  wire                ifm_sign_x_1_14;
  wire                ifm_sign_x_1_15;
  wire                ifm_sign_x_1_16;
  wire                ifm_sign_x_2_0;
  wire                ifm_sign_x_2_1;
  wire                ifm_sign_x_2_2;
  wire                ifm_sign_x_2_3;
  wire                ifm_sign_x_2_4;
  wire                ifm_sign_x_2_5;
  wire                ifm_sign_x_2_6;
  wire                ifm_sign_x_2_7;
  wire                ifm_sign_x_2_8;
  wire                ifm_sign_x_2_9;
  wire                ifm_sign_x_2_10;
  wire                ifm_sign_x_2_11;
  wire                ifm_sign_x_2_12;
  wire                ifm_sign_x_2_13;
  wire                ifm_sign_x_2_14;
  wire                ifm_sign_x_2_15;
  wire                ifm_sign_x_2_16;
  wire                ifm_sign_x_3_0;
  wire                ifm_sign_x_3_1;
  wire                ifm_sign_x_3_2;
  wire                ifm_sign_x_3_3;
  wire                ifm_sign_x_3_4;
  wire                ifm_sign_x_3_5;
  wire                ifm_sign_x_3_6;
  wire                ifm_sign_x_3_7;
  wire                ifm_sign_x_3_8;
  wire                ifm_sign_x_3_9;
  wire                ifm_sign_x_3_10;
  wire                ifm_sign_x_3_11;
  wire                ifm_sign_x_3_12;
  wire                ifm_sign_x_3_13;
  wire                ifm_sign_x_3_14;
  wire                ifm_sign_x_3_15;
  wire                ifm_sign_x_3_16;
  wire                ifm_sign_x_4_0;
  wire                ifm_sign_x_4_1;
  wire                ifm_sign_x_4_2;
  wire                ifm_sign_x_4_3;
  wire                ifm_sign_x_4_4;
  wire                ifm_sign_x_4_5;
  wire                ifm_sign_x_4_6;
  wire                ifm_sign_x_4_7;
  wire                ifm_sign_x_4_8;
  wire                ifm_sign_x_4_9;
  wire                ifm_sign_x_4_10;
  wire                ifm_sign_x_4_11;
  wire                ifm_sign_x_4_12;
  wire                ifm_sign_x_4_13;
  wire                ifm_sign_x_4_14;
  wire                ifm_sign_x_4_15;
  wire                ifm_sign_x_4_16;
  wire                ifm_sign_x_5_0;
  wire                ifm_sign_x_5_1;
  wire                ifm_sign_x_5_2;
  wire                ifm_sign_x_5_3;
  wire                ifm_sign_x_5_4;
  wire                ifm_sign_x_5_5;
  wire                ifm_sign_x_5_6;
  wire                ifm_sign_x_5_7;
  wire                ifm_sign_x_5_8;
  wire                ifm_sign_x_5_9;
  wire                ifm_sign_x_5_10;
  wire                ifm_sign_x_5_11;
  wire                ifm_sign_x_5_12;
  wire                ifm_sign_x_5_13;
  wire                ifm_sign_x_5_14;
  wire                ifm_sign_x_5_15;
  wire                ifm_sign_x_5_16;
  wire                ifm_sign_x_6_0;
  wire                ifm_sign_x_6_1;
  wire                ifm_sign_x_6_2;
  wire                ifm_sign_x_6_3;
  wire                ifm_sign_x_6_4;
  wire                ifm_sign_x_6_5;
  wire                ifm_sign_x_6_6;
  wire                ifm_sign_x_6_7;
  wire                ifm_sign_x_6_8;
  wire                ifm_sign_x_6_9;
  wire                ifm_sign_x_6_10;
  wire                ifm_sign_x_6_11;
  wire                ifm_sign_x_6_12;
  wire                ifm_sign_x_6_13;
  wire                ifm_sign_x_6_14;
  wire                ifm_sign_x_6_15;
  wire                ifm_sign_x_6_16;
  wire                ifm_sign_x_7_0;
  wire                ifm_sign_x_7_1;
  wire                ifm_sign_x_7_2;
  wire                ifm_sign_x_7_3;
  wire                ifm_sign_x_7_4;
  wire                ifm_sign_x_7_5;
  wire                ifm_sign_x_7_6;
  wire                ifm_sign_x_7_7;
  wire                ifm_sign_x_7_8;
  wire                ifm_sign_x_7_9;
  wire                ifm_sign_x_7_10;
  wire                ifm_sign_x_7_11;
  wire                ifm_sign_x_7_12;
  wire                ifm_sign_x_7_13;
  wire                ifm_sign_x_7_14;
  wire                ifm_sign_x_7_15;
  wire                ifm_sign_x_7_16;
  wire                ifm_sign_x_8_0;
  wire                ifm_sign_x_8_1;
  wire                ifm_sign_x_8_2;
  wire                ifm_sign_x_8_3;
  wire                ifm_sign_x_8_4;
  wire                ifm_sign_x_8_5;
  wire                ifm_sign_x_8_6;
  wire                ifm_sign_x_8_7;
  wire                ifm_sign_x_8_8;
  wire                ifm_sign_x_8_9;
  wire                ifm_sign_x_8_10;
  wire                ifm_sign_x_8_11;
  wire                ifm_sign_x_8_12;
  wire                ifm_sign_x_8_13;
  wire                ifm_sign_x_8_14;
  wire                ifm_sign_x_8_15;
  wire                ifm_sign_x_8_16;
  wire                ifm_sign_x_9_0;
  wire                ifm_sign_x_9_1;
  wire                ifm_sign_x_9_2;
  wire                ifm_sign_x_9_3;
  wire                ifm_sign_x_9_4;
  wire                ifm_sign_x_9_5;
  wire                ifm_sign_x_9_6;
  wire                ifm_sign_x_9_7;
  wire                ifm_sign_x_9_8;
  wire                ifm_sign_x_9_9;
  wire                ifm_sign_x_9_10;
  wire                ifm_sign_x_9_11;
  wire                ifm_sign_x_9_12;
  wire                ifm_sign_x_9_13;
  wire                ifm_sign_x_9_14;
  wire                ifm_sign_x_9_15;
  wire                ifm_sign_x_9_16;
  wire                ifm_sign_x_10_0;
  wire                ifm_sign_x_10_1;
  wire                ifm_sign_x_10_2;
  wire                ifm_sign_x_10_3;
  wire                ifm_sign_x_10_4;
  wire                ifm_sign_x_10_5;
  wire                ifm_sign_x_10_6;
  wire                ifm_sign_x_10_7;
  wire                ifm_sign_x_10_8;
  wire                ifm_sign_x_10_9;
  wire                ifm_sign_x_10_10;
  wire                ifm_sign_x_10_11;
  wire                ifm_sign_x_10_12;
  wire                ifm_sign_x_10_13;
  wire                ifm_sign_x_10_14;
  wire                ifm_sign_x_10_15;
  wire                ifm_sign_x_10_16;
  wire                ifm_sign_x_11_0;
  wire                ifm_sign_x_11_1;
  wire                ifm_sign_x_11_2;
  wire                ifm_sign_x_11_3;
  wire                ifm_sign_x_11_4;
  wire                ifm_sign_x_11_5;
  wire                ifm_sign_x_11_6;
  wire                ifm_sign_x_11_7;
  wire                ifm_sign_x_11_8;
  wire                ifm_sign_x_11_9;
  wire                ifm_sign_x_11_10;
  wire                ifm_sign_x_11_11;
  wire                ifm_sign_x_11_12;
  wire                ifm_sign_x_11_13;
  wire                ifm_sign_x_11_14;
  wire                ifm_sign_x_11_15;
  wire                ifm_sign_x_11_16;
  wire                ifm_sign_x_12_0;
  wire                ifm_sign_x_12_1;
  wire                ifm_sign_x_12_2;
  wire                ifm_sign_x_12_3;
  wire                ifm_sign_x_12_4;
  wire                ifm_sign_x_12_5;
  wire                ifm_sign_x_12_6;
  wire                ifm_sign_x_12_7;
  wire                ifm_sign_x_12_8;
  wire                ifm_sign_x_12_9;
  wire                ifm_sign_x_12_10;
  wire                ifm_sign_x_12_11;
  wire                ifm_sign_x_12_12;
  wire                ifm_sign_x_12_13;
  wire                ifm_sign_x_12_14;
  wire                ifm_sign_x_12_15;
  wire                ifm_sign_x_12_16;
  wire                ifm_sign_x_13_0;
  wire                ifm_sign_x_13_1;
  wire                ifm_sign_x_13_2;
  wire                ifm_sign_x_13_3;
  wire                ifm_sign_x_13_4;
  wire                ifm_sign_x_13_5;
  wire                ifm_sign_x_13_6;
  wire                ifm_sign_x_13_7;
  wire                ifm_sign_x_13_8;
  wire                ifm_sign_x_13_9;
  wire                ifm_sign_x_13_10;
  wire                ifm_sign_x_13_11;
  wire                ifm_sign_x_13_12;
  wire                ifm_sign_x_13_13;
  wire                ifm_sign_x_13_14;
  wire                ifm_sign_x_13_15;
  wire                ifm_sign_x_13_16;
  wire                ifm_sign_x_14_0;
  wire                ifm_sign_x_14_1;
  wire                ifm_sign_x_14_2;
  wire                ifm_sign_x_14_3;
  wire                ifm_sign_x_14_4;
  wire                ifm_sign_x_14_5;
  wire                ifm_sign_x_14_6;
  wire                ifm_sign_x_14_7;
  wire                ifm_sign_x_14_8;
  wire                ifm_sign_x_14_9;
  wire                ifm_sign_x_14_10;
  wire                ifm_sign_x_14_11;
  wire                ifm_sign_x_14_12;
  wire                ifm_sign_x_14_13;
  wire                ifm_sign_x_14_14;
  wire                ifm_sign_x_14_15;
  wire                ifm_sign_x_14_16;
  wire                ifm_sign_x_15_0;
  wire                ifm_sign_x_15_1;
  wire                ifm_sign_x_15_2;
  wire                ifm_sign_x_15_3;
  wire                ifm_sign_x_15_4;
  wire                ifm_sign_x_15_5;
  wire                ifm_sign_x_15_6;
  wire                ifm_sign_x_15_7;
  wire                ifm_sign_x_15_8;
  wire                ifm_sign_x_15_9;
  wire                ifm_sign_x_15_10;
  wire                ifm_sign_x_15_11;
  wire                ifm_sign_x_15_12;
  wire                ifm_sign_x_15_13;
  wire                ifm_sign_x_15_14;
  wire                ifm_sign_x_15_15;
  wire                ifm_sign_x_15_16;
  wire                ifm_dff_x_0_0;
  wire                ifm_dff_x_0_1;
  wire                ifm_dff_x_0_2;
  wire                ifm_dff_x_0_3;
  wire                ifm_dff_x_0_4;
  wire                ifm_dff_x_0_5;
  wire                ifm_dff_x_0_6;
  wire                ifm_dff_x_0_7;
  wire                ifm_dff_x_0_8;
  wire                ifm_dff_x_0_9;
  wire                ifm_dff_x_0_10;
  wire                ifm_dff_x_0_11;
  wire                ifm_dff_x_0_12;
  wire                ifm_dff_x_0_13;
  wire                ifm_dff_x_0_14;
  wire                ifm_dff_x_0_15;
  wire                ifm_dff_x_0_16;
  wire                ifm_dff_x_1_0;
  wire                ifm_dff_x_1_1;
  wire                ifm_dff_x_1_2;
  wire                ifm_dff_x_1_3;
  wire                ifm_dff_x_1_4;
  wire                ifm_dff_x_1_5;
  wire                ifm_dff_x_1_6;
  wire                ifm_dff_x_1_7;
  wire                ifm_dff_x_1_8;
  wire                ifm_dff_x_1_9;
  wire                ifm_dff_x_1_10;
  wire                ifm_dff_x_1_11;
  wire                ifm_dff_x_1_12;
  wire                ifm_dff_x_1_13;
  wire                ifm_dff_x_1_14;
  wire                ifm_dff_x_1_15;
  wire                ifm_dff_x_1_16;
  wire                ifm_dff_x_2_0;
  wire                ifm_dff_x_2_1;
  wire                ifm_dff_x_2_2;
  wire                ifm_dff_x_2_3;
  wire                ifm_dff_x_2_4;
  wire                ifm_dff_x_2_5;
  wire                ifm_dff_x_2_6;
  wire                ifm_dff_x_2_7;
  wire                ifm_dff_x_2_8;
  wire                ifm_dff_x_2_9;
  wire                ifm_dff_x_2_10;
  wire                ifm_dff_x_2_11;
  wire                ifm_dff_x_2_12;
  wire                ifm_dff_x_2_13;
  wire                ifm_dff_x_2_14;
  wire                ifm_dff_x_2_15;
  wire                ifm_dff_x_2_16;
  wire                ifm_dff_x_3_0;
  wire                ifm_dff_x_3_1;
  wire                ifm_dff_x_3_2;
  wire                ifm_dff_x_3_3;
  wire                ifm_dff_x_3_4;
  wire                ifm_dff_x_3_5;
  wire                ifm_dff_x_3_6;
  wire                ifm_dff_x_3_7;
  wire                ifm_dff_x_3_8;
  wire                ifm_dff_x_3_9;
  wire                ifm_dff_x_3_10;
  wire                ifm_dff_x_3_11;
  wire                ifm_dff_x_3_12;
  wire                ifm_dff_x_3_13;
  wire                ifm_dff_x_3_14;
  wire                ifm_dff_x_3_15;
  wire                ifm_dff_x_3_16;
  wire                ifm_dff_x_4_0;
  wire                ifm_dff_x_4_1;
  wire                ifm_dff_x_4_2;
  wire                ifm_dff_x_4_3;
  wire                ifm_dff_x_4_4;
  wire                ifm_dff_x_4_5;
  wire                ifm_dff_x_4_6;
  wire                ifm_dff_x_4_7;
  wire                ifm_dff_x_4_8;
  wire                ifm_dff_x_4_9;
  wire                ifm_dff_x_4_10;
  wire                ifm_dff_x_4_11;
  wire                ifm_dff_x_4_12;
  wire                ifm_dff_x_4_13;
  wire                ifm_dff_x_4_14;
  wire                ifm_dff_x_4_15;
  wire                ifm_dff_x_4_16;
  wire                ifm_dff_x_5_0;
  wire                ifm_dff_x_5_1;
  wire                ifm_dff_x_5_2;
  wire                ifm_dff_x_5_3;
  wire                ifm_dff_x_5_4;
  wire                ifm_dff_x_5_5;
  wire                ifm_dff_x_5_6;
  wire                ifm_dff_x_5_7;
  wire                ifm_dff_x_5_8;
  wire                ifm_dff_x_5_9;
  wire                ifm_dff_x_5_10;
  wire                ifm_dff_x_5_11;
  wire                ifm_dff_x_5_12;
  wire                ifm_dff_x_5_13;
  wire                ifm_dff_x_5_14;
  wire                ifm_dff_x_5_15;
  wire                ifm_dff_x_5_16;
  wire                ifm_dff_x_6_0;
  wire                ifm_dff_x_6_1;
  wire                ifm_dff_x_6_2;
  wire                ifm_dff_x_6_3;
  wire                ifm_dff_x_6_4;
  wire                ifm_dff_x_6_5;
  wire                ifm_dff_x_6_6;
  wire                ifm_dff_x_6_7;
  wire                ifm_dff_x_6_8;
  wire                ifm_dff_x_6_9;
  wire                ifm_dff_x_6_10;
  wire                ifm_dff_x_6_11;
  wire                ifm_dff_x_6_12;
  wire                ifm_dff_x_6_13;
  wire                ifm_dff_x_6_14;
  wire                ifm_dff_x_6_15;
  wire                ifm_dff_x_6_16;
  wire                ifm_dff_x_7_0;
  wire                ifm_dff_x_7_1;
  wire                ifm_dff_x_7_2;
  wire                ifm_dff_x_7_3;
  wire                ifm_dff_x_7_4;
  wire                ifm_dff_x_7_5;
  wire                ifm_dff_x_7_6;
  wire                ifm_dff_x_7_7;
  wire                ifm_dff_x_7_8;
  wire                ifm_dff_x_7_9;
  wire                ifm_dff_x_7_10;
  wire                ifm_dff_x_7_11;
  wire                ifm_dff_x_7_12;
  wire                ifm_dff_x_7_13;
  wire                ifm_dff_x_7_14;
  wire                ifm_dff_x_7_15;
  wire                ifm_dff_x_7_16;
  wire                ifm_dff_x_8_0;
  wire                ifm_dff_x_8_1;
  wire                ifm_dff_x_8_2;
  wire                ifm_dff_x_8_3;
  wire                ifm_dff_x_8_4;
  wire                ifm_dff_x_8_5;
  wire                ifm_dff_x_8_6;
  wire                ifm_dff_x_8_7;
  wire                ifm_dff_x_8_8;
  wire                ifm_dff_x_8_9;
  wire                ifm_dff_x_8_10;
  wire                ifm_dff_x_8_11;
  wire                ifm_dff_x_8_12;
  wire                ifm_dff_x_8_13;
  wire                ifm_dff_x_8_14;
  wire                ifm_dff_x_8_15;
  wire                ifm_dff_x_8_16;
  wire                ifm_dff_x_9_0;
  wire                ifm_dff_x_9_1;
  wire                ifm_dff_x_9_2;
  wire                ifm_dff_x_9_3;
  wire                ifm_dff_x_9_4;
  wire                ifm_dff_x_9_5;
  wire                ifm_dff_x_9_6;
  wire                ifm_dff_x_9_7;
  wire                ifm_dff_x_9_8;
  wire                ifm_dff_x_9_9;
  wire                ifm_dff_x_9_10;
  wire                ifm_dff_x_9_11;
  wire                ifm_dff_x_9_12;
  wire                ifm_dff_x_9_13;
  wire                ifm_dff_x_9_14;
  wire                ifm_dff_x_9_15;
  wire                ifm_dff_x_9_16;
  wire                ifm_dff_x_10_0;
  wire                ifm_dff_x_10_1;
  wire                ifm_dff_x_10_2;
  wire                ifm_dff_x_10_3;
  wire                ifm_dff_x_10_4;
  wire                ifm_dff_x_10_5;
  wire                ifm_dff_x_10_6;
  wire                ifm_dff_x_10_7;
  wire                ifm_dff_x_10_8;
  wire                ifm_dff_x_10_9;
  wire                ifm_dff_x_10_10;
  wire                ifm_dff_x_10_11;
  wire                ifm_dff_x_10_12;
  wire                ifm_dff_x_10_13;
  wire                ifm_dff_x_10_14;
  wire                ifm_dff_x_10_15;
  wire                ifm_dff_x_10_16;
  wire                ifm_dff_x_11_0;
  wire                ifm_dff_x_11_1;
  wire                ifm_dff_x_11_2;
  wire                ifm_dff_x_11_3;
  wire                ifm_dff_x_11_4;
  wire                ifm_dff_x_11_5;
  wire                ifm_dff_x_11_6;
  wire                ifm_dff_x_11_7;
  wire                ifm_dff_x_11_8;
  wire                ifm_dff_x_11_9;
  wire                ifm_dff_x_11_10;
  wire                ifm_dff_x_11_11;
  wire                ifm_dff_x_11_12;
  wire                ifm_dff_x_11_13;
  wire                ifm_dff_x_11_14;
  wire                ifm_dff_x_11_15;
  wire                ifm_dff_x_11_16;
  wire                ifm_dff_x_12_0;
  wire                ifm_dff_x_12_1;
  wire                ifm_dff_x_12_2;
  wire                ifm_dff_x_12_3;
  wire                ifm_dff_x_12_4;
  wire                ifm_dff_x_12_5;
  wire                ifm_dff_x_12_6;
  wire                ifm_dff_x_12_7;
  wire                ifm_dff_x_12_8;
  wire                ifm_dff_x_12_9;
  wire                ifm_dff_x_12_10;
  wire                ifm_dff_x_12_11;
  wire                ifm_dff_x_12_12;
  wire                ifm_dff_x_12_13;
  wire                ifm_dff_x_12_14;
  wire                ifm_dff_x_12_15;
  wire                ifm_dff_x_12_16;
  wire                ifm_dff_x_13_0;
  wire                ifm_dff_x_13_1;
  wire                ifm_dff_x_13_2;
  wire                ifm_dff_x_13_3;
  wire                ifm_dff_x_13_4;
  wire                ifm_dff_x_13_5;
  wire                ifm_dff_x_13_6;
  wire                ifm_dff_x_13_7;
  wire                ifm_dff_x_13_8;
  wire                ifm_dff_x_13_9;
  wire                ifm_dff_x_13_10;
  wire                ifm_dff_x_13_11;
  wire                ifm_dff_x_13_12;
  wire                ifm_dff_x_13_13;
  wire                ifm_dff_x_13_14;
  wire                ifm_dff_x_13_15;
  wire                ifm_dff_x_13_16;
  wire                ifm_dff_x_14_0;
  wire                ifm_dff_x_14_1;
  wire                ifm_dff_x_14_2;
  wire                ifm_dff_x_14_3;
  wire                ifm_dff_x_14_4;
  wire                ifm_dff_x_14_5;
  wire                ifm_dff_x_14_6;
  wire                ifm_dff_x_14_7;
  wire                ifm_dff_x_14_8;
  wire                ifm_dff_x_14_9;
  wire                ifm_dff_x_14_10;
  wire                ifm_dff_x_14_11;
  wire                ifm_dff_x_14_12;
  wire                ifm_dff_x_14_13;
  wire                ifm_dff_x_14_14;
  wire                ifm_dff_x_14_15;
  wire                ifm_dff_x_14_16;
  wire                ifm_dff_x_15_0;
  wire                ifm_dff_x_15_1;
  wire                ifm_dff_x_15_2;
  wire                ifm_dff_x_15_3;
  wire                ifm_dff_x_15_4;
  wire                ifm_dff_x_15_5;
  wire                ifm_dff_x_15_6;
  wire                ifm_dff_x_15_7;
  wire                ifm_dff_x_15_8;
  wire                ifm_dff_x_15_9;
  wire                ifm_dff_x_15_10;
  wire                ifm_dff_x_15_11;
  wire                ifm_dff_x_15_12;
  wire                ifm_dff_x_15_13;
  wire                ifm_dff_x_15_14;
  wire                ifm_dff_x_15_15;
  wire                ifm_dff_x_15_16;
  wire                wght_sign_x_0_0;
  wire                wght_sign_x_0_1;
  wire                wght_sign_x_0_2;
  wire                wght_sign_x_0_3;
  wire                wght_sign_x_0_4;
  wire                wght_sign_x_0_5;
  wire                wght_sign_x_0_6;
  wire                wght_sign_x_0_7;
  wire                wght_sign_x_0_8;
  wire                wght_sign_x_0_9;
  wire                wght_sign_x_0_10;
  wire                wght_sign_x_0_11;
  wire                wght_sign_x_0_12;
  wire                wght_sign_x_0_13;
  wire                wght_sign_x_0_14;
  wire                wght_sign_x_0_15;
  wire                wght_sign_x_0_16;
  wire                wght_sign_x_1_0;
  wire                wght_sign_x_1_1;
  wire                wght_sign_x_1_2;
  wire                wght_sign_x_1_3;
  wire                wght_sign_x_1_4;
  wire                wght_sign_x_1_5;
  wire                wght_sign_x_1_6;
  wire                wght_sign_x_1_7;
  wire                wght_sign_x_1_8;
  wire                wght_sign_x_1_9;
  wire                wght_sign_x_1_10;
  wire                wght_sign_x_1_11;
  wire                wght_sign_x_1_12;
  wire                wght_sign_x_1_13;
  wire                wght_sign_x_1_14;
  wire                wght_sign_x_1_15;
  wire                wght_sign_x_1_16;
  wire                wght_sign_x_2_0;
  wire                wght_sign_x_2_1;
  wire                wght_sign_x_2_2;
  wire                wght_sign_x_2_3;
  wire                wght_sign_x_2_4;
  wire                wght_sign_x_2_5;
  wire                wght_sign_x_2_6;
  wire                wght_sign_x_2_7;
  wire                wght_sign_x_2_8;
  wire                wght_sign_x_2_9;
  wire                wght_sign_x_2_10;
  wire                wght_sign_x_2_11;
  wire                wght_sign_x_2_12;
  wire                wght_sign_x_2_13;
  wire                wght_sign_x_2_14;
  wire                wght_sign_x_2_15;
  wire                wght_sign_x_2_16;
  wire                wght_sign_x_3_0;
  wire                wght_sign_x_3_1;
  wire                wght_sign_x_3_2;
  wire                wght_sign_x_3_3;
  wire                wght_sign_x_3_4;
  wire                wght_sign_x_3_5;
  wire                wght_sign_x_3_6;
  wire                wght_sign_x_3_7;
  wire                wght_sign_x_3_8;
  wire                wght_sign_x_3_9;
  wire                wght_sign_x_3_10;
  wire                wght_sign_x_3_11;
  wire                wght_sign_x_3_12;
  wire                wght_sign_x_3_13;
  wire                wght_sign_x_3_14;
  wire                wght_sign_x_3_15;
  wire                wght_sign_x_3_16;
  wire                wght_sign_x_4_0;
  wire                wght_sign_x_4_1;
  wire                wght_sign_x_4_2;
  wire                wght_sign_x_4_3;
  wire                wght_sign_x_4_4;
  wire                wght_sign_x_4_5;
  wire                wght_sign_x_4_6;
  wire                wght_sign_x_4_7;
  wire                wght_sign_x_4_8;
  wire                wght_sign_x_4_9;
  wire                wght_sign_x_4_10;
  wire                wght_sign_x_4_11;
  wire                wght_sign_x_4_12;
  wire                wght_sign_x_4_13;
  wire                wght_sign_x_4_14;
  wire                wght_sign_x_4_15;
  wire                wght_sign_x_4_16;
  wire                wght_sign_x_5_0;
  wire                wght_sign_x_5_1;
  wire                wght_sign_x_5_2;
  wire                wght_sign_x_5_3;
  wire                wght_sign_x_5_4;
  wire                wght_sign_x_5_5;
  wire                wght_sign_x_5_6;
  wire                wght_sign_x_5_7;
  wire                wght_sign_x_5_8;
  wire                wght_sign_x_5_9;
  wire                wght_sign_x_5_10;
  wire                wght_sign_x_5_11;
  wire                wght_sign_x_5_12;
  wire                wght_sign_x_5_13;
  wire                wght_sign_x_5_14;
  wire                wght_sign_x_5_15;
  wire                wght_sign_x_5_16;
  wire                wght_sign_x_6_0;
  wire                wght_sign_x_6_1;
  wire                wght_sign_x_6_2;
  wire                wght_sign_x_6_3;
  wire                wght_sign_x_6_4;
  wire                wght_sign_x_6_5;
  wire                wght_sign_x_6_6;
  wire                wght_sign_x_6_7;
  wire                wght_sign_x_6_8;
  wire                wght_sign_x_6_9;
  wire                wght_sign_x_6_10;
  wire                wght_sign_x_6_11;
  wire                wght_sign_x_6_12;
  wire                wght_sign_x_6_13;
  wire                wght_sign_x_6_14;
  wire                wght_sign_x_6_15;
  wire                wght_sign_x_6_16;
  wire                wght_sign_x_7_0;
  wire                wght_sign_x_7_1;
  wire                wght_sign_x_7_2;
  wire                wght_sign_x_7_3;
  wire                wght_sign_x_7_4;
  wire                wght_sign_x_7_5;
  wire                wght_sign_x_7_6;
  wire                wght_sign_x_7_7;
  wire                wght_sign_x_7_8;
  wire                wght_sign_x_7_9;
  wire                wght_sign_x_7_10;
  wire                wght_sign_x_7_11;
  wire                wght_sign_x_7_12;
  wire                wght_sign_x_7_13;
  wire                wght_sign_x_7_14;
  wire                wght_sign_x_7_15;
  wire                wght_sign_x_7_16;
  wire                wght_sign_x_8_0;
  wire                wght_sign_x_8_1;
  wire                wght_sign_x_8_2;
  wire                wght_sign_x_8_3;
  wire                wght_sign_x_8_4;
  wire                wght_sign_x_8_5;
  wire                wght_sign_x_8_6;
  wire                wght_sign_x_8_7;
  wire                wght_sign_x_8_8;
  wire                wght_sign_x_8_9;
  wire                wght_sign_x_8_10;
  wire                wght_sign_x_8_11;
  wire                wght_sign_x_8_12;
  wire                wght_sign_x_8_13;
  wire                wght_sign_x_8_14;
  wire                wght_sign_x_8_15;
  wire                wght_sign_x_8_16;
  wire                wght_sign_x_9_0;
  wire                wght_sign_x_9_1;
  wire                wght_sign_x_9_2;
  wire                wght_sign_x_9_3;
  wire                wght_sign_x_9_4;
  wire                wght_sign_x_9_5;
  wire                wght_sign_x_9_6;
  wire                wght_sign_x_9_7;
  wire                wght_sign_x_9_8;
  wire                wght_sign_x_9_9;
  wire                wght_sign_x_9_10;
  wire                wght_sign_x_9_11;
  wire                wght_sign_x_9_12;
  wire                wght_sign_x_9_13;
  wire                wght_sign_x_9_14;
  wire                wght_sign_x_9_15;
  wire                wght_sign_x_9_16;
  wire                wght_sign_x_10_0;
  wire                wght_sign_x_10_1;
  wire                wght_sign_x_10_2;
  wire                wght_sign_x_10_3;
  wire                wght_sign_x_10_4;
  wire                wght_sign_x_10_5;
  wire                wght_sign_x_10_6;
  wire                wght_sign_x_10_7;
  wire                wght_sign_x_10_8;
  wire                wght_sign_x_10_9;
  wire                wght_sign_x_10_10;
  wire                wght_sign_x_10_11;
  wire                wght_sign_x_10_12;
  wire                wght_sign_x_10_13;
  wire                wght_sign_x_10_14;
  wire                wght_sign_x_10_15;
  wire                wght_sign_x_10_16;
  wire                wght_sign_x_11_0;
  wire                wght_sign_x_11_1;
  wire                wght_sign_x_11_2;
  wire                wght_sign_x_11_3;
  wire                wght_sign_x_11_4;
  wire                wght_sign_x_11_5;
  wire                wght_sign_x_11_6;
  wire                wght_sign_x_11_7;
  wire                wght_sign_x_11_8;
  wire                wght_sign_x_11_9;
  wire                wght_sign_x_11_10;
  wire                wght_sign_x_11_11;
  wire                wght_sign_x_11_12;
  wire                wght_sign_x_11_13;
  wire                wght_sign_x_11_14;
  wire                wght_sign_x_11_15;
  wire                wght_sign_x_11_16;
  wire                wght_sign_x_12_0;
  wire                wght_sign_x_12_1;
  wire                wght_sign_x_12_2;
  wire                wght_sign_x_12_3;
  wire                wght_sign_x_12_4;
  wire                wght_sign_x_12_5;
  wire                wght_sign_x_12_6;
  wire                wght_sign_x_12_7;
  wire                wght_sign_x_12_8;
  wire                wght_sign_x_12_9;
  wire                wght_sign_x_12_10;
  wire                wght_sign_x_12_11;
  wire                wght_sign_x_12_12;
  wire                wght_sign_x_12_13;
  wire                wght_sign_x_12_14;
  wire                wght_sign_x_12_15;
  wire                wght_sign_x_12_16;
  wire                wght_sign_x_13_0;
  wire                wght_sign_x_13_1;
  wire                wght_sign_x_13_2;
  wire                wght_sign_x_13_3;
  wire                wght_sign_x_13_4;
  wire                wght_sign_x_13_5;
  wire                wght_sign_x_13_6;
  wire                wght_sign_x_13_7;
  wire                wght_sign_x_13_8;
  wire                wght_sign_x_13_9;
  wire                wght_sign_x_13_10;
  wire                wght_sign_x_13_11;
  wire                wght_sign_x_13_12;
  wire                wght_sign_x_13_13;
  wire                wght_sign_x_13_14;
  wire                wght_sign_x_13_15;
  wire                wght_sign_x_13_16;
  wire                wght_sign_x_14_0;
  wire                wght_sign_x_14_1;
  wire                wght_sign_x_14_2;
  wire                wght_sign_x_14_3;
  wire                wght_sign_x_14_4;
  wire                wght_sign_x_14_5;
  wire                wght_sign_x_14_6;
  wire                wght_sign_x_14_7;
  wire                wght_sign_x_14_8;
  wire                wght_sign_x_14_9;
  wire                wght_sign_x_14_10;
  wire                wght_sign_x_14_11;
  wire                wght_sign_x_14_12;
  wire                wght_sign_x_14_13;
  wire                wght_sign_x_14_14;
  wire                wght_sign_x_14_15;
  wire                wght_sign_x_14_16;
  wire                wght_sign_x_15_0;
  wire                wght_sign_x_15_1;
  wire                wght_sign_x_15_2;
  wire                wght_sign_x_15_3;
  wire                wght_sign_x_15_4;
  wire                wght_sign_x_15_5;
  wire                wght_sign_x_15_6;
  wire                wght_sign_x_15_7;
  wire                wght_sign_x_15_8;
  wire                wght_sign_x_15_9;
  wire                wght_sign_x_15_10;
  wire                wght_sign_x_15_11;
  wire                wght_sign_x_15_12;
  wire                wght_sign_x_15_13;
  wire                wght_sign_x_15_14;
  wire                wght_sign_x_15_15;
  wire                wght_sign_x_15_16;
  wire       [14:0]   wght_abs_x_0_0;
  wire       [14:0]   wght_abs_x_0_1;
  wire       [14:0]   wght_abs_x_0_2;
  wire       [14:0]   wght_abs_x_0_3;
  wire       [14:0]   wght_abs_x_0_4;
  wire       [14:0]   wght_abs_x_0_5;
  wire       [14:0]   wght_abs_x_0_6;
  wire       [14:0]   wght_abs_x_0_7;
  wire       [14:0]   wght_abs_x_0_8;
  wire       [14:0]   wght_abs_x_0_9;
  wire       [14:0]   wght_abs_x_0_10;
  wire       [14:0]   wght_abs_x_0_11;
  wire       [14:0]   wght_abs_x_0_12;
  wire       [14:0]   wght_abs_x_0_13;
  wire       [14:0]   wght_abs_x_0_14;
  wire       [14:0]   wght_abs_x_0_15;
  wire       [14:0]   wght_abs_x_0_16;
  wire       [14:0]   wght_abs_x_1_0;
  wire       [14:0]   wght_abs_x_1_1;
  wire       [14:0]   wght_abs_x_1_2;
  wire       [14:0]   wght_abs_x_1_3;
  wire       [14:0]   wght_abs_x_1_4;
  wire       [14:0]   wght_abs_x_1_5;
  wire       [14:0]   wght_abs_x_1_6;
  wire       [14:0]   wght_abs_x_1_7;
  wire       [14:0]   wght_abs_x_1_8;
  wire       [14:0]   wght_abs_x_1_9;
  wire       [14:0]   wght_abs_x_1_10;
  wire       [14:0]   wght_abs_x_1_11;
  wire       [14:0]   wght_abs_x_1_12;
  wire       [14:0]   wght_abs_x_1_13;
  wire       [14:0]   wght_abs_x_1_14;
  wire       [14:0]   wght_abs_x_1_15;
  wire       [14:0]   wght_abs_x_1_16;
  wire       [14:0]   wght_abs_x_2_0;
  wire       [14:0]   wght_abs_x_2_1;
  wire       [14:0]   wght_abs_x_2_2;
  wire       [14:0]   wght_abs_x_2_3;
  wire       [14:0]   wght_abs_x_2_4;
  wire       [14:0]   wght_abs_x_2_5;
  wire       [14:0]   wght_abs_x_2_6;
  wire       [14:0]   wght_abs_x_2_7;
  wire       [14:0]   wght_abs_x_2_8;
  wire       [14:0]   wght_abs_x_2_9;
  wire       [14:0]   wght_abs_x_2_10;
  wire       [14:0]   wght_abs_x_2_11;
  wire       [14:0]   wght_abs_x_2_12;
  wire       [14:0]   wght_abs_x_2_13;
  wire       [14:0]   wght_abs_x_2_14;
  wire       [14:0]   wght_abs_x_2_15;
  wire       [14:0]   wght_abs_x_2_16;
  wire       [14:0]   wght_abs_x_3_0;
  wire       [14:0]   wght_abs_x_3_1;
  wire       [14:0]   wght_abs_x_3_2;
  wire       [14:0]   wght_abs_x_3_3;
  wire       [14:0]   wght_abs_x_3_4;
  wire       [14:0]   wght_abs_x_3_5;
  wire       [14:0]   wght_abs_x_3_6;
  wire       [14:0]   wght_abs_x_3_7;
  wire       [14:0]   wght_abs_x_3_8;
  wire       [14:0]   wght_abs_x_3_9;
  wire       [14:0]   wght_abs_x_3_10;
  wire       [14:0]   wght_abs_x_3_11;
  wire       [14:0]   wght_abs_x_3_12;
  wire       [14:0]   wght_abs_x_3_13;
  wire       [14:0]   wght_abs_x_3_14;
  wire       [14:0]   wght_abs_x_3_15;
  wire       [14:0]   wght_abs_x_3_16;
  wire       [14:0]   wght_abs_x_4_0;
  wire       [14:0]   wght_abs_x_4_1;
  wire       [14:0]   wght_abs_x_4_2;
  wire       [14:0]   wght_abs_x_4_3;
  wire       [14:0]   wght_abs_x_4_4;
  wire       [14:0]   wght_abs_x_4_5;
  wire       [14:0]   wght_abs_x_4_6;
  wire       [14:0]   wght_abs_x_4_7;
  wire       [14:0]   wght_abs_x_4_8;
  wire       [14:0]   wght_abs_x_4_9;
  wire       [14:0]   wght_abs_x_4_10;
  wire       [14:0]   wght_abs_x_4_11;
  wire       [14:0]   wght_abs_x_4_12;
  wire       [14:0]   wght_abs_x_4_13;
  wire       [14:0]   wght_abs_x_4_14;
  wire       [14:0]   wght_abs_x_4_15;
  wire       [14:0]   wght_abs_x_4_16;
  wire       [14:0]   wght_abs_x_5_0;
  wire       [14:0]   wght_abs_x_5_1;
  wire       [14:0]   wght_abs_x_5_2;
  wire       [14:0]   wght_abs_x_5_3;
  wire       [14:0]   wght_abs_x_5_4;
  wire       [14:0]   wght_abs_x_5_5;
  wire       [14:0]   wght_abs_x_5_6;
  wire       [14:0]   wght_abs_x_5_7;
  wire       [14:0]   wght_abs_x_5_8;
  wire       [14:0]   wght_abs_x_5_9;
  wire       [14:0]   wght_abs_x_5_10;
  wire       [14:0]   wght_abs_x_5_11;
  wire       [14:0]   wght_abs_x_5_12;
  wire       [14:0]   wght_abs_x_5_13;
  wire       [14:0]   wght_abs_x_5_14;
  wire       [14:0]   wght_abs_x_5_15;
  wire       [14:0]   wght_abs_x_5_16;
  wire       [14:0]   wght_abs_x_6_0;
  wire       [14:0]   wght_abs_x_6_1;
  wire       [14:0]   wght_abs_x_6_2;
  wire       [14:0]   wght_abs_x_6_3;
  wire       [14:0]   wght_abs_x_6_4;
  wire       [14:0]   wght_abs_x_6_5;
  wire       [14:0]   wght_abs_x_6_6;
  wire       [14:0]   wght_abs_x_6_7;
  wire       [14:0]   wght_abs_x_6_8;
  wire       [14:0]   wght_abs_x_6_9;
  wire       [14:0]   wght_abs_x_6_10;
  wire       [14:0]   wght_abs_x_6_11;
  wire       [14:0]   wght_abs_x_6_12;
  wire       [14:0]   wght_abs_x_6_13;
  wire       [14:0]   wght_abs_x_6_14;
  wire       [14:0]   wght_abs_x_6_15;
  wire       [14:0]   wght_abs_x_6_16;
  wire       [14:0]   wght_abs_x_7_0;
  wire       [14:0]   wght_abs_x_7_1;
  wire       [14:0]   wght_abs_x_7_2;
  wire       [14:0]   wght_abs_x_7_3;
  wire       [14:0]   wght_abs_x_7_4;
  wire       [14:0]   wght_abs_x_7_5;
  wire       [14:0]   wght_abs_x_7_6;
  wire       [14:0]   wght_abs_x_7_7;
  wire       [14:0]   wght_abs_x_7_8;
  wire       [14:0]   wght_abs_x_7_9;
  wire       [14:0]   wght_abs_x_7_10;
  wire       [14:0]   wght_abs_x_7_11;
  wire       [14:0]   wght_abs_x_7_12;
  wire       [14:0]   wght_abs_x_7_13;
  wire       [14:0]   wght_abs_x_7_14;
  wire       [14:0]   wght_abs_x_7_15;
  wire       [14:0]   wght_abs_x_7_16;
  wire       [14:0]   wght_abs_x_8_0;
  wire       [14:0]   wght_abs_x_8_1;
  wire       [14:0]   wght_abs_x_8_2;
  wire       [14:0]   wght_abs_x_8_3;
  wire       [14:0]   wght_abs_x_8_4;
  wire       [14:0]   wght_abs_x_8_5;
  wire       [14:0]   wght_abs_x_8_6;
  wire       [14:0]   wght_abs_x_8_7;
  wire       [14:0]   wght_abs_x_8_8;
  wire       [14:0]   wght_abs_x_8_9;
  wire       [14:0]   wght_abs_x_8_10;
  wire       [14:0]   wght_abs_x_8_11;
  wire       [14:0]   wght_abs_x_8_12;
  wire       [14:0]   wght_abs_x_8_13;
  wire       [14:0]   wght_abs_x_8_14;
  wire       [14:0]   wght_abs_x_8_15;
  wire       [14:0]   wght_abs_x_8_16;
  wire       [14:0]   wght_abs_x_9_0;
  wire       [14:0]   wght_abs_x_9_1;
  wire       [14:0]   wght_abs_x_9_2;
  wire       [14:0]   wght_abs_x_9_3;
  wire       [14:0]   wght_abs_x_9_4;
  wire       [14:0]   wght_abs_x_9_5;
  wire       [14:0]   wght_abs_x_9_6;
  wire       [14:0]   wght_abs_x_9_7;
  wire       [14:0]   wght_abs_x_9_8;
  wire       [14:0]   wght_abs_x_9_9;
  wire       [14:0]   wght_abs_x_9_10;
  wire       [14:0]   wght_abs_x_9_11;
  wire       [14:0]   wght_abs_x_9_12;
  wire       [14:0]   wght_abs_x_9_13;
  wire       [14:0]   wght_abs_x_9_14;
  wire       [14:0]   wght_abs_x_9_15;
  wire       [14:0]   wght_abs_x_9_16;
  wire       [14:0]   wght_abs_x_10_0;
  wire       [14:0]   wght_abs_x_10_1;
  wire       [14:0]   wght_abs_x_10_2;
  wire       [14:0]   wght_abs_x_10_3;
  wire       [14:0]   wght_abs_x_10_4;
  wire       [14:0]   wght_abs_x_10_5;
  wire       [14:0]   wght_abs_x_10_6;
  wire       [14:0]   wght_abs_x_10_7;
  wire       [14:0]   wght_abs_x_10_8;
  wire       [14:0]   wght_abs_x_10_9;
  wire       [14:0]   wght_abs_x_10_10;
  wire       [14:0]   wght_abs_x_10_11;
  wire       [14:0]   wght_abs_x_10_12;
  wire       [14:0]   wght_abs_x_10_13;
  wire       [14:0]   wght_abs_x_10_14;
  wire       [14:0]   wght_abs_x_10_15;
  wire       [14:0]   wght_abs_x_10_16;
  wire       [14:0]   wght_abs_x_11_0;
  wire       [14:0]   wght_abs_x_11_1;
  wire       [14:0]   wght_abs_x_11_2;
  wire       [14:0]   wght_abs_x_11_3;
  wire       [14:0]   wght_abs_x_11_4;
  wire       [14:0]   wght_abs_x_11_5;
  wire       [14:0]   wght_abs_x_11_6;
  wire       [14:0]   wght_abs_x_11_7;
  wire       [14:0]   wght_abs_x_11_8;
  wire       [14:0]   wght_abs_x_11_9;
  wire       [14:0]   wght_abs_x_11_10;
  wire       [14:0]   wght_abs_x_11_11;
  wire       [14:0]   wght_abs_x_11_12;
  wire       [14:0]   wght_abs_x_11_13;
  wire       [14:0]   wght_abs_x_11_14;
  wire       [14:0]   wght_abs_x_11_15;
  wire       [14:0]   wght_abs_x_11_16;
  wire       [14:0]   wght_abs_x_12_0;
  wire       [14:0]   wght_abs_x_12_1;
  wire       [14:0]   wght_abs_x_12_2;
  wire       [14:0]   wght_abs_x_12_3;
  wire       [14:0]   wght_abs_x_12_4;
  wire       [14:0]   wght_abs_x_12_5;
  wire       [14:0]   wght_abs_x_12_6;
  wire       [14:0]   wght_abs_x_12_7;
  wire       [14:0]   wght_abs_x_12_8;
  wire       [14:0]   wght_abs_x_12_9;
  wire       [14:0]   wght_abs_x_12_10;
  wire       [14:0]   wght_abs_x_12_11;
  wire       [14:0]   wght_abs_x_12_12;
  wire       [14:0]   wght_abs_x_12_13;
  wire       [14:0]   wght_abs_x_12_14;
  wire       [14:0]   wght_abs_x_12_15;
  wire       [14:0]   wght_abs_x_12_16;
  wire       [14:0]   wght_abs_x_13_0;
  wire       [14:0]   wght_abs_x_13_1;
  wire       [14:0]   wght_abs_x_13_2;
  wire       [14:0]   wght_abs_x_13_3;
  wire       [14:0]   wght_abs_x_13_4;
  wire       [14:0]   wght_abs_x_13_5;
  wire       [14:0]   wght_abs_x_13_6;
  wire       [14:0]   wght_abs_x_13_7;
  wire       [14:0]   wght_abs_x_13_8;
  wire       [14:0]   wght_abs_x_13_9;
  wire       [14:0]   wght_abs_x_13_10;
  wire       [14:0]   wght_abs_x_13_11;
  wire       [14:0]   wght_abs_x_13_12;
  wire       [14:0]   wght_abs_x_13_13;
  wire       [14:0]   wght_abs_x_13_14;
  wire       [14:0]   wght_abs_x_13_15;
  wire       [14:0]   wght_abs_x_13_16;
  wire       [14:0]   wght_abs_x_14_0;
  wire       [14:0]   wght_abs_x_14_1;
  wire       [14:0]   wght_abs_x_14_2;
  wire       [14:0]   wght_abs_x_14_3;
  wire       [14:0]   wght_abs_x_14_4;
  wire       [14:0]   wght_abs_x_14_5;
  wire       [14:0]   wght_abs_x_14_6;
  wire       [14:0]   wght_abs_x_14_7;
  wire       [14:0]   wght_abs_x_14_8;
  wire       [14:0]   wght_abs_x_14_9;
  wire       [14:0]   wght_abs_x_14_10;
  wire       [14:0]   wght_abs_x_14_11;
  wire       [14:0]   wght_abs_x_14_12;
  wire       [14:0]   wght_abs_x_14_13;
  wire       [14:0]   wght_abs_x_14_14;
  wire       [14:0]   wght_abs_x_14_15;
  wire       [14:0]   wght_abs_x_14_16;
  wire       [14:0]   wght_abs_x_15_0;
  wire       [14:0]   wght_abs_x_15_1;
  wire       [14:0]   wght_abs_x_15_2;
  wire       [14:0]   wght_abs_x_15_3;
  wire       [14:0]   wght_abs_x_15_4;
  wire       [14:0]   wght_abs_x_15_5;
  wire       [14:0]   wght_abs_x_15_6;
  wire       [14:0]   wght_abs_x_15_7;
  wire       [14:0]   wght_abs_x_15_8;
  wire       [14:0]   wght_abs_x_15_9;
  wire       [14:0]   wght_abs_x_15_10;
  wire       [14:0]   wght_abs_x_15_11;
  wire       [14:0]   wght_abs_x_15_12;
  wire       [14:0]   wght_abs_x_15_13;
  wire       [14:0]   wght_abs_x_15_14;
  wire       [14:0]   wght_abs_x_15_15;
  wire       [14:0]   wght_abs_x_15_16;
  wire       [14:0]   randW_x_0_0;
  wire       [14:0]   randW_x_0_1;
  wire       [14:0]   randW_x_0_2;
  wire       [14:0]   randW_x_0_3;
  wire       [14:0]   randW_x_0_4;
  wire       [14:0]   randW_x_0_5;
  wire       [14:0]   randW_x_0_6;
  wire       [14:0]   randW_x_0_7;
  wire       [14:0]   randW_x_0_8;
  wire       [14:0]   randW_x_0_9;
  wire       [14:0]   randW_x_0_10;
  wire       [14:0]   randW_x_0_11;
  wire       [14:0]   randW_x_0_12;
  wire       [14:0]   randW_x_0_13;
  wire       [14:0]   randW_x_0_14;
  wire       [14:0]   randW_x_0_15;
  wire       [14:0]   randW_x_0_16;
  wire       [14:0]   randW_x_1_0;
  wire       [14:0]   randW_x_1_1;
  wire       [14:0]   randW_x_1_2;
  wire       [14:0]   randW_x_1_3;
  wire       [14:0]   randW_x_1_4;
  wire       [14:0]   randW_x_1_5;
  wire       [14:0]   randW_x_1_6;
  wire       [14:0]   randW_x_1_7;
  wire       [14:0]   randW_x_1_8;
  wire       [14:0]   randW_x_1_9;
  wire       [14:0]   randW_x_1_10;
  wire       [14:0]   randW_x_1_11;
  wire       [14:0]   randW_x_1_12;
  wire       [14:0]   randW_x_1_13;
  wire       [14:0]   randW_x_1_14;
  wire       [14:0]   randW_x_1_15;
  wire       [14:0]   randW_x_1_16;
  wire       [14:0]   randW_x_2_0;
  wire       [14:0]   randW_x_2_1;
  wire       [14:0]   randW_x_2_2;
  wire       [14:0]   randW_x_2_3;
  wire       [14:0]   randW_x_2_4;
  wire       [14:0]   randW_x_2_5;
  wire       [14:0]   randW_x_2_6;
  wire       [14:0]   randW_x_2_7;
  wire       [14:0]   randW_x_2_8;
  wire       [14:0]   randW_x_2_9;
  wire       [14:0]   randW_x_2_10;
  wire       [14:0]   randW_x_2_11;
  wire       [14:0]   randW_x_2_12;
  wire       [14:0]   randW_x_2_13;
  wire       [14:0]   randW_x_2_14;
  wire       [14:0]   randW_x_2_15;
  wire       [14:0]   randW_x_2_16;
  wire       [14:0]   randW_x_3_0;
  wire       [14:0]   randW_x_3_1;
  wire       [14:0]   randW_x_3_2;
  wire       [14:0]   randW_x_3_3;
  wire       [14:0]   randW_x_3_4;
  wire       [14:0]   randW_x_3_5;
  wire       [14:0]   randW_x_3_6;
  wire       [14:0]   randW_x_3_7;
  wire       [14:0]   randW_x_3_8;
  wire       [14:0]   randW_x_3_9;
  wire       [14:0]   randW_x_3_10;
  wire       [14:0]   randW_x_3_11;
  wire       [14:0]   randW_x_3_12;
  wire       [14:0]   randW_x_3_13;
  wire       [14:0]   randW_x_3_14;
  wire       [14:0]   randW_x_3_15;
  wire       [14:0]   randW_x_3_16;
  wire       [14:0]   randW_x_4_0;
  wire       [14:0]   randW_x_4_1;
  wire       [14:0]   randW_x_4_2;
  wire       [14:0]   randW_x_4_3;
  wire       [14:0]   randW_x_4_4;
  wire       [14:0]   randW_x_4_5;
  wire       [14:0]   randW_x_4_6;
  wire       [14:0]   randW_x_4_7;
  wire       [14:0]   randW_x_4_8;
  wire       [14:0]   randW_x_4_9;
  wire       [14:0]   randW_x_4_10;
  wire       [14:0]   randW_x_4_11;
  wire       [14:0]   randW_x_4_12;
  wire       [14:0]   randW_x_4_13;
  wire       [14:0]   randW_x_4_14;
  wire       [14:0]   randW_x_4_15;
  wire       [14:0]   randW_x_4_16;
  wire       [14:0]   randW_x_5_0;
  wire       [14:0]   randW_x_5_1;
  wire       [14:0]   randW_x_5_2;
  wire       [14:0]   randW_x_5_3;
  wire       [14:0]   randW_x_5_4;
  wire       [14:0]   randW_x_5_5;
  wire       [14:0]   randW_x_5_6;
  wire       [14:0]   randW_x_5_7;
  wire       [14:0]   randW_x_5_8;
  wire       [14:0]   randW_x_5_9;
  wire       [14:0]   randW_x_5_10;
  wire       [14:0]   randW_x_5_11;
  wire       [14:0]   randW_x_5_12;
  wire       [14:0]   randW_x_5_13;
  wire       [14:0]   randW_x_5_14;
  wire       [14:0]   randW_x_5_15;
  wire       [14:0]   randW_x_5_16;
  wire       [14:0]   randW_x_6_0;
  wire       [14:0]   randW_x_6_1;
  wire       [14:0]   randW_x_6_2;
  wire       [14:0]   randW_x_6_3;
  wire       [14:0]   randW_x_6_4;
  wire       [14:0]   randW_x_6_5;
  wire       [14:0]   randW_x_6_6;
  wire       [14:0]   randW_x_6_7;
  wire       [14:0]   randW_x_6_8;
  wire       [14:0]   randW_x_6_9;
  wire       [14:0]   randW_x_6_10;
  wire       [14:0]   randW_x_6_11;
  wire       [14:0]   randW_x_6_12;
  wire       [14:0]   randW_x_6_13;
  wire       [14:0]   randW_x_6_14;
  wire       [14:0]   randW_x_6_15;
  wire       [14:0]   randW_x_6_16;
  wire       [14:0]   randW_x_7_0;
  wire       [14:0]   randW_x_7_1;
  wire       [14:0]   randW_x_7_2;
  wire       [14:0]   randW_x_7_3;
  wire       [14:0]   randW_x_7_4;
  wire       [14:0]   randW_x_7_5;
  wire       [14:0]   randW_x_7_6;
  wire       [14:0]   randW_x_7_7;
  wire       [14:0]   randW_x_7_8;
  wire       [14:0]   randW_x_7_9;
  wire       [14:0]   randW_x_7_10;
  wire       [14:0]   randW_x_7_11;
  wire       [14:0]   randW_x_7_12;
  wire       [14:0]   randW_x_7_13;
  wire       [14:0]   randW_x_7_14;
  wire       [14:0]   randW_x_7_15;
  wire       [14:0]   randW_x_7_16;
  wire       [14:0]   randW_x_8_0;
  wire       [14:0]   randW_x_8_1;
  wire       [14:0]   randW_x_8_2;
  wire       [14:0]   randW_x_8_3;
  wire       [14:0]   randW_x_8_4;
  wire       [14:0]   randW_x_8_5;
  wire       [14:0]   randW_x_8_6;
  wire       [14:0]   randW_x_8_7;
  wire       [14:0]   randW_x_8_8;
  wire       [14:0]   randW_x_8_9;
  wire       [14:0]   randW_x_8_10;
  wire       [14:0]   randW_x_8_11;
  wire       [14:0]   randW_x_8_12;
  wire       [14:0]   randW_x_8_13;
  wire       [14:0]   randW_x_8_14;
  wire       [14:0]   randW_x_8_15;
  wire       [14:0]   randW_x_8_16;
  wire       [14:0]   randW_x_9_0;
  wire       [14:0]   randW_x_9_1;
  wire       [14:0]   randW_x_9_2;
  wire       [14:0]   randW_x_9_3;
  wire       [14:0]   randW_x_9_4;
  wire       [14:0]   randW_x_9_5;
  wire       [14:0]   randW_x_9_6;
  wire       [14:0]   randW_x_9_7;
  wire       [14:0]   randW_x_9_8;
  wire       [14:0]   randW_x_9_9;
  wire       [14:0]   randW_x_9_10;
  wire       [14:0]   randW_x_9_11;
  wire       [14:0]   randW_x_9_12;
  wire       [14:0]   randW_x_9_13;
  wire       [14:0]   randW_x_9_14;
  wire       [14:0]   randW_x_9_15;
  wire       [14:0]   randW_x_9_16;
  wire       [14:0]   randW_x_10_0;
  wire       [14:0]   randW_x_10_1;
  wire       [14:0]   randW_x_10_2;
  wire       [14:0]   randW_x_10_3;
  wire       [14:0]   randW_x_10_4;
  wire       [14:0]   randW_x_10_5;
  wire       [14:0]   randW_x_10_6;
  wire       [14:0]   randW_x_10_7;
  wire       [14:0]   randW_x_10_8;
  wire       [14:0]   randW_x_10_9;
  wire       [14:0]   randW_x_10_10;
  wire       [14:0]   randW_x_10_11;
  wire       [14:0]   randW_x_10_12;
  wire       [14:0]   randW_x_10_13;
  wire       [14:0]   randW_x_10_14;
  wire       [14:0]   randW_x_10_15;
  wire       [14:0]   randW_x_10_16;
  wire       [14:0]   randW_x_11_0;
  wire       [14:0]   randW_x_11_1;
  wire       [14:0]   randW_x_11_2;
  wire       [14:0]   randW_x_11_3;
  wire       [14:0]   randW_x_11_4;
  wire       [14:0]   randW_x_11_5;
  wire       [14:0]   randW_x_11_6;
  wire       [14:0]   randW_x_11_7;
  wire       [14:0]   randW_x_11_8;
  wire       [14:0]   randW_x_11_9;
  wire       [14:0]   randW_x_11_10;
  wire       [14:0]   randW_x_11_11;
  wire       [14:0]   randW_x_11_12;
  wire       [14:0]   randW_x_11_13;
  wire       [14:0]   randW_x_11_14;
  wire       [14:0]   randW_x_11_15;
  wire       [14:0]   randW_x_11_16;
  wire       [14:0]   randW_x_12_0;
  wire       [14:0]   randW_x_12_1;
  wire       [14:0]   randW_x_12_2;
  wire       [14:0]   randW_x_12_3;
  wire       [14:0]   randW_x_12_4;
  wire       [14:0]   randW_x_12_5;
  wire       [14:0]   randW_x_12_6;
  wire       [14:0]   randW_x_12_7;
  wire       [14:0]   randW_x_12_8;
  wire       [14:0]   randW_x_12_9;
  wire       [14:0]   randW_x_12_10;
  wire       [14:0]   randW_x_12_11;
  wire       [14:0]   randW_x_12_12;
  wire       [14:0]   randW_x_12_13;
  wire       [14:0]   randW_x_12_14;
  wire       [14:0]   randW_x_12_15;
  wire       [14:0]   randW_x_12_16;
  wire       [14:0]   randW_x_13_0;
  wire       [14:0]   randW_x_13_1;
  wire       [14:0]   randW_x_13_2;
  wire       [14:0]   randW_x_13_3;
  wire       [14:0]   randW_x_13_4;
  wire       [14:0]   randW_x_13_5;
  wire       [14:0]   randW_x_13_6;
  wire       [14:0]   randW_x_13_7;
  wire       [14:0]   randW_x_13_8;
  wire       [14:0]   randW_x_13_9;
  wire       [14:0]   randW_x_13_10;
  wire       [14:0]   randW_x_13_11;
  wire       [14:0]   randW_x_13_12;
  wire       [14:0]   randW_x_13_13;
  wire       [14:0]   randW_x_13_14;
  wire       [14:0]   randW_x_13_15;
  wire       [14:0]   randW_x_13_16;
  wire       [14:0]   randW_x_14_0;
  wire       [14:0]   randW_x_14_1;
  wire       [14:0]   randW_x_14_2;
  wire       [14:0]   randW_x_14_3;
  wire       [14:0]   randW_x_14_4;
  wire       [14:0]   randW_x_14_5;
  wire       [14:0]   randW_x_14_6;
  wire       [14:0]   randW_x_14_7;
  wire       [14:0]   randW_x_14_8;
  wire       [14:0]   randW_x_14_9;
  wire       [14:0]   randW_x_14_10;
  wire       [14:0]   randW_x_14_11;
  wire       [14:0]   randW_x_14_12;
  wire       [14:0]   randW_x_14_13;
  wire       [14:0]   randW_x_14_14;
  wire       [14:0]   randW_x_14_15;
  wire       [14:0]   randW_x_14_16;
  wire       [14:0]   randW_x_15_0;
  wire       [14:0]   randW_x_15_1;
  wire       [14:0]   randW_x_15_2;
  wire       [14:0]   randW_x_15_3;
  wire       [14:0]   randW_x_15_4;
  wire       [14:0]   randW_x_15_5;
  wire       [14:0]   randW_x_15_6;
  wire       [14:0]   randW_x_15_7;
  wire       [14:0]   randW_x_15_8;
  wire       [14:0]   randW_x_15_9;
  wire       [14:0]   randW_x_15_10;
  wire       [14:0]   randW_x_15_11;
  wire       [14:0]   randW_x_15_12;
  wire       [14:0]   randW_x_15_13;
  wire       [14:0]   randW_x_15_14;
  wire       [14:0]   randW_x_15_15;
  wire       [14:0]   randW_x_15_16;
  wire       [31:0]   ofm_x_0_0;
  wire       [31:0]   ofm_x_0_1;
  wire       [31:0]   ofm_x_0_2;
  wire       [31:0]   ofm_x_0_3;
  wire       [31:0]   ofm_x_0_4;
  wire       [31:0]   ofm_x_0_5;
  wire       [31:0]   ofm_x_0_6;
  wire       [31:0]   ofm_x_0_7;
  wire       [31:0]   ofm_x_0_8;
  wire       [31:0]   ofm_x_0_9;
  wire       [31:0]   ofm_x_0_10;
  wire       [31:0]   ofm_x_0_11;
  wire       [31:0]   ofm_x_0_12;
  wire       [31:0]   ofm_x_0_13;
  wire       [31:0]   ofm_x_0_14;
  wire       [31:0]   ofm_x_0_15;
  wire       [31:0]   ofm_x_0_16;
  wire       [31:0]   ofm_x_1_0;
  wire       [31:0]   ofm_x_1_1;
  wire       [31:0]   ofm_x_1_2;
  wire       [31:0]   ofm_x_1_3;
  wire       [31:0]   ofm_x_1_4;
  wire       [31:0]   ofm_x_1_5;
  wire       [31:0]   ofm_x_1_6;
  wire       [31:0]   ofm_x_1_7;
  wire       [31:0]   ofm_x_1_8;
  wire       [31:0]   ofm_x_1_9;
  wire       [31:0]   ofm_x_1_10;
  wire       [31:0]   ofm_x_1_11;
  wire       [31:0]   ofm_x_1_12;
  wire       [31:0]   ofm_x_1_13;
  wire       [31:0]   ofm_x_1_14;
  wire       [31:0]   ofm_x_1_15;
  wire       [31:0]   ofm_x_1_16;
  wire       [31:0]   ofm_x_2_0;
  wire       [31:0]   ofm_x_2_1;
  wire       [31:0]   ofm_x_2_2;
  wire       [31:0]   ofm_x_2_3;
  wire       [31:0]   ofm_x_2_4;
  wire       [31:0]   ofm_x_2_5;
  wire       [31:0]   ofm_x_2_6;
  wire       [31:0]   ofm_x_2_7;
  wire       [31:0]   ofm_x_2_8;
  wire       [31:0]   ofm_x_2_9;
  wire       [31:0]   ofm_x_2_10;
  wire       [31:0]   ofm_x_2_11;
  wire       [31:0]   ofm_x_2_12;
  wire       [31:0]   ofm_x_2_13;
  wire       [31:0]   ofm_x_2_14;
  wire       [31:0]   ofm_x_2_15;
  wire       [31:0]   ofm_x_2_16;
  wire       [31:0]   ofm_x_3_0;
  wire       [31:0]   ofm_x_3_1;
  wire       [31:0]   ofm_x_3_2;
  wire       [31:0]   ofm_x_3_3;
  wire       [31:0]   ofm_x_3_4;
  wire       [31:0]   ofm_x_3_5;
  wire       [31:0]   ofm_x_3_6;
  wire       [31:0]   ofm_x_3_7;
  wire       [31:0]   ofm_x_3_8;
  wire       [31:0]   ofm_x_3_9;
  wire       [31:0]   ofm_x_3_10;
  wire       [31:0]   ofm_x_3_11;
  wire       [31:0]   ofm_x_3_12;
  wire       [31:0]   ofm_x_3_13;
  wire       [31:0]   ofm_x_3_14;
  wire       [31:0]   ofm_x_3_15;
  wire       [31:0]   ofm_x_3_16;
  wire       [31:0]   ofm_x_4_0;
  wire       [31:0]   ofm_x_4_1;
  wire       [31:0]   ofm_x_4_2;
  wire       [31:0]   ofm_x_4_3;
  wire       [31:0]   ofm_x_4_4;
  wire       [31:0]   ofm_x_4_5;
  wire       [31:0]   ofm_x_4_6;
  wire       [31:0]   ofm_x_4_7;
  wire       [31:0]   ofm_x_4_8;
  wire       [31:0]   ofm_x_4_9;
  wire       [31:0]   ofm_x_4_10;
  wire       [31:0]   ofm_x_4_11;
  wire       [31:0]   ofm_x_4_12;
  wire       [31:0]   ofm_x_4_13;
  wire       [31:0]   ofm_x_4_14;
  wire       [31:0]   ofm_x_4_15;
  wire       [31:0]   ofm_x_4_16;
  wire       [31:0]   ofm_x_5_0;
  wire       [31:0]   ofm_x_5_1;
  wire       [31:0]   ofm_x_5_2;
  wire       [31:0]   ofm_x_5_3;
  wire       [31:0]   ofm_x_5_4;
  wire       [31:0]   ofm_x_5_5;
  wire       [31:0]   ofm_x_5_6;
  wire       [31:0]   ofm_x_5_7;
  wire       [31:0]   ofm_x_5_8;
  wire       [31:0]   ofm_x_5_9;
  wire       [31:0]   ofm_x_5_10;
  wire       [31:0]   ofm_x_5_11;
  wire       [31:0]   ofm_x_5_12;
  wire       [31:0]   ofm_x_5_13;
  wire       [31:0]   ofm_x_5_14;
  wire       [31:0]   ofm_x_5_15;
  wire       [31:0]   ofm_x_5_16;
  wire       [31:0]   ofm_x_6_0;
  wire       [31:0]   ofm_x_6_1;
  wire       [31:0]   ofm_x_6_2;
  wire       [31:0]   ofm_x_6_3;
  wire       [31:0]   ofm_x_6_4;
  wire       [31:0]   ofm_x_6_5;
  wire       [31:0]   ofm_x_6_6;
  wire       [31:0]   ofm_x_6_7;
  wire       [31:0]   ofm_x_6_8;
  wire       [31:0]   ofm_x_6_9;
  wire       [31:0]   ofm_x_6_10;
  wire       [31:0]   ofm_x_6_11;
  wire       [31:0]   ofm_x_6_12;
  wire       [31:0]   ofm_x_6_13;
  wire       [31:0]   ofm_x_6_14;
  wire       [31:0]   ofm_x_6_15;
  wire       [31:0]   ofm_x_6_16;
  wire       [31:0]   ofm_x_7_0;
  wire       [31:0]   ofm_x_7_1;
  wire       [31:0]   ofm_x_7_2;
  wire       [31:0]   ofm_x_7_3;
  wire       [31:0]   ofm_x_7_4;
  wire       [31:0]   ofm_x_7_5;
  wire       [31:0]   ofm_x_7_6;
  wire       [31:0]   ofm_x_7_7;
  wire       [31:0]   ofm_x_7_8;
  wire       [31:0]   ofm_x_7_9;
  wire       [31:0]   ofm_x_7_10;
  wire       [31:0]   ofm_x_7_11;
  wire       [31:0]   ofm_x_7_12;
  wire       [31:0]   ofm_x_7_13;
  wire       [31:0]   ofm_x_7_14;
  wire       [31:0]   ofm_x_7_15;
  wire       [31:0]   ofm_x_7_16;
  wire       [31:0]   ofm_x_8_0;
  wire       [31:0]   ofm_x_8_1;
  wire       [31:0]   ofm_x_8_2;
  wire       [31:0]   ofm_x_8_3;
  wire       [31:0]   ofm_x_8_4;
  wire       [31:0]   ofm_x_8_5;
  wire       [31:0]   ofm_x_8_6;
  wire       [31:0]   ofm_x_8_7;
  wire       [31:0]   ofm_x_8_8;
  wire       [31:0]   ofm_x_8_9;
  wire       [31:0]   ofm_x_8_10;
  wire       [31:0]   ofm_x_8_11;
  wire       [31:0]   ofm_x_8_12;
  wire       [31:0]   ofm_x_8_13;
  wire       [31:0]   ofm_x_8_14;
  wire       [31:0]   ofm_x_8_15;
  wire       [31:0]   ofm_x_8_16;
  wire       [31:0]   ofm_x_9_0;
  wire       [31:0]   ofm_x_9_1;
  wire       [31:0]   ofm_x_9_2;
  wire       [31:0]   ofm_x_9_3;
  wire       [31:0]   ofm_x_9_4;
  wire       [31:0]   ofm_x_9_5;
  wire       [31:0]   ofm_x_9_6;
  wire       [31:0]   ofm_x_9_7;
  wire       [31:0]   ofm_x_9_8;
  wire       [31:0]   ofm_x_9_9;
  wire       [31:0]   ofm_x_9_10;
  wire       [31:0]   ofm_x_9_11;
  wire       [31:0]   ofm_x_9_12;
  wire       [31:0]   ofm_x_9_13;
  wire       [31:0]   ofm_x_9_14;
  wire       [31:0]   ofm_x_9_15;
  wire       [31:0]   ofm_x_9_16;
  wire       [31:0]   ofm_x_10_0;
  wire       [31:0]   ofm_x_10_1;
  wire       [31:0]   ofm_x_10_2;
  wire       [31:0]   ofm_x_10_3;
  wire       [31:0]   ofm_x_10_4;
  wire       [31:0]   ofm_x_10_5;
  wire       [31:0]   ofm_x_10_6;
  wire       [31:0]   ofm_x_10_7;
  wire       [31:0]   ofm_x_10_8;
  wire       [31:0]   ofm_x_10_9;
  wire       [31:0]   ofm_x_10_10;
  wire       [31:0]   ofm_x_10_11;
  wire       [31:0]   ofm_x_10_12;
  wire       [31:0]   ofm_x_10_13;
  wire       [31:0]   ofm_x_10_14;
  wire       [31:0]   ofm_x_10_15;
  wire       [31:0]   ofm_x_10_16;
  wire       [31:0]   ofm_x_11_0;
  wire       [31:0]   ofm_x_11_1;
  wire       [31:0]   ofm_x_11_2;
  wire       [31:0]   ofm_x_11_3;
  wire       [31:0]   ofm_x_11_4;
  wire       [31:0]   ofm_x_11_5;
  wire       [31:0]   ofm_x_11_6;
  wire       [31:0]   ofm_x_11_7;
  wire       [31:0]   ofm_x_11_8;
  wire       [31:0]   ofm_x_11_9;
  wire       [31:0]   ofm_x_11_10;
  wire       [31:0]   ofm_x_11_11;
  wire       [31:0]   ofm_x_11_12;
  wire       [31:0]   ofm_x_11_13;
  wire       [31:0]   ofm_x_11_14;
  wire       [31:0]   ofm_x_11_15;
  wire       [31:0]   ofm_x_11_16;
  wire       [31:0]   ofm_x_12_0;
  wire       [31:0]   ofm_x_12_1;
  wire       [31:0]   ofm_x_12_2;
  wire       [31:0]   ofm_x_12_3;
  wire       [31:0]   ofm_x_12_4;
  wire       [31:0]   ofm_x_12_5;
  wire       [31:0]   ofm_x_12_6;
  wire       [31:0]   ofm_x_12_7;
  wire       [31:0]   ofm_x_12_8;
  wire       [31:0]   ofm_x_12_9;
  wire       [31:0]   ofm_x_12_10;
  wire       [31:0]   ofm_x_12_11;
  wire       [31:0]   ofm_x_12_12;
  wire       [31:0]   ofm_x_12_13;
  wire       [31:0]   ofm_x_12_14;
  wire       [31:0]   ofm_x_12_15;
  wire       [31:0]   ofm_x_12_16;
  wire       [31:0]   ofm_x_13_0;
  wire       [31:0]   ofm_x_13_1;
  wire       [31:0]   ofm_x_13_2;
  wire       [31:0]   ofm_x_13_3;
  wire       [31:0]   ofm_x_13_4;
  wire       [31:0]   ofm_x_13_5;
  wire       [31:0]   ofm_x_13_6;
  wire       [31:0]   ofm_x_13_7;
  wire       [31:0]   ofm_x_13_8;
  wire       [31:0]   ofm_x_13_9;
  wire       [31:0]   ofm_x_13_10;
  wire       [31:0]   ofm_x_13_11;
  wire       [31:0]   ofm_x_13_12;
  wire       [31:0]   ofm_x_13_13;
  wire       [31:0]   ofm_x_13_14;
  wire       [31:0]   ofm_x_13_15;
  wire       [31:0]   ofm_x_13_16;
  wire       [31:0]   ofm_x_14_0;
  wire       [31:0]   ofm_x_14_1;
  wire       [31:0]   ofm_x_14_2;
  wire       [31:0]   ofm_x_14_3;
  wire       [31:0]   ofm_x_14_4;
  wire       [31:0]   ofm_x_14_5;
  wire       [31:0]   ofm_x_14_6;
  wire       [31:0]   ofm_x_14_7;
  wire       [31:0]   ofm_x_14_8;
  wire       [31:0]   ofm_x_14_9;
  wire       [31:0]   ofm_x_14_10;
  wire       [31:0]   ofm_x_14_11;
  wire       [31:0]   ofm_x_14_12;
  wire       [31:0]   ofm_x_14_13;
  wire       [31:0]   ofm_x_14_14;
  wire       [31:0]   ofm_x_14_15;
  wire       [31:0]   ofm_x_14_16;
  wire       [31:0]   ofm_x_15_0;
  wire       [31:0]   ofm_x_15_1;
  wire       [31:0]   ofm_x_15_2;
  wire       [31:0]   ofm_x_15_3;
  wire       [31:0]   ofm_x_15_4;
  wire       [31:0]   ofm_x_15_5;
  wire       [31:0]   ofm_x_15_6;
  wire       [31:0]   ofm_x_15_7;
  wire       [31:0]   ofm_x_15_8;
  wire       [31:0]   ofm_x_15_9;
  wire       [31:0]   ofm_x_15_10;
  wire       [31:0]   ofm_x_15_11;
  wire       [31:0]   ofm_x_15_12;
  wire       [31:0]   ofm_x_15_13;
  wire       [31:0]   ofm_x_15_14;
  wire       [31:0]   ofm_x_15_15;
  wire       [31:0]   ofm_x_15_16;

  uSystolicPEBorder uSystolicPEBorder_16 (
    .io_mac_done    (uSystolicPEBorder_16_io_mac_done        ), //i
    .io_enable_i    (uSystolicPEBorder_16_io_enable_i        ), //i
    .io_clear_i     (uSystolicPEBorder_16_io_clear_i         ), //i
    .io_enable_w    (uSystolicPEBorder_16_io_enable_w        ), //i
    .io_clear_w     (uSystolicPEBorder_16_io_clear_w         ), //i
    .io_enable_o    (uSystolicPEBorder_16_io_enable_o        ), //i
    .io_clear_o     (uSystolicPEBorder_16_io_clear_o         ), //i
    .io_ifm         (io_ifm_0[15:0]                          ), //i
    .io_wght_sign   (wght_sign_x_0_0                         ), //i
    .io_wght_abs    (wght_abs_x_0_0[14:0]                    ), //i
    .io_ofm         (ofm_x_0_1[31:0]                         ), //i
    .io_mac_done_d  (uSystolicPEBorder_16_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPEBorder_16_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPEBorder_16_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPEBorder_16_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPEBorder_16_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPEBorder_16_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPEBorder_16_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPEBorder_16_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPEBorder_16_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPEBorder_16_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPEBorder_16_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPEBorder_16_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPEBorder_16_io_ofm_d[31:0]     ), //o
    .clk            (clk                                     ), //i
    .reset          (reset                                   )  //i
  );
  uSystolicPE uSystolicPE_240 (
    .io_mac_done    (uSystolicPE_240_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_240_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_240_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_240_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_240_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_240_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_240_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_0_1                     ), //i
    .io_ifm_dff     (ifm_dff_x_0_1                      ), //i
    .io_wght_sign   (wght_sign_x_1_0                    ), //i
    .io_randW       (randW_x_0_1[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_1_0[14:0]               ), //i
    .io_ofm         (ofm_x_1_1[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_240_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_240_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_240_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_240_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_240_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_240_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_240_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_240_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_240_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_240_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_240_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_240_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_240_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_241 (
    .io_mac_done    (uSystolicPE_241_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_241_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_241_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_241_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_241_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_241_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_241_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_0_2                     ), //i
    .io_ifm_dff     (ifm_dff_x_0_2                      ), //i
    .io_wght_sign   (wght_sign_x_2_0                    ), //i
    .io_randW       (randW_x_0_2[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_2_0[14:0]               ), //i
    .io_ofm         (ofm_x_2_1[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_241_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_241_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_241_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_241_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_241_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_241_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_241_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_241_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_241_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_241_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_241_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_241_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_241_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_242 (
    .io_mac_done    (uSystolicPE_242_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_242_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_242_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_242_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_242_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_242_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_242_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_0_3                     ), //i
    .io_ifm_dff     (ifm_dff_x_0_3                      ), //i
    .io_wght_sign   (wght_sign_x_3_0                    ), //i
    .io_randW       (randW_x_0_3[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_3_0[14:0]               ), //i
    .io_ofm         (ofm_x_3_1[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_242_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_242_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_242_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_242_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_242_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_242_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_242_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_242_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_242_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_242_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_242_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_242_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_242_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_243 (
    .io_mac_done    (uSystolicPE_243_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_243_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_243_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_243_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_243_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_243_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_243_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_0_4                     ), //i
    .io_ifm_dff     (ifm_dff_x_0_4                      ), //i
    .io_wght_sign   (wght_sign_x_4_0                    ), //i
    .io_randW       (randW_x_0_4[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_4_0[14:0]               ), //i
    .io_ofm         (ofm_x_4_1[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_243_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_243_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_243_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_243_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_243_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_243_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_243_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_243_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_243_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_243_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_243_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_243_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_243_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_244 (
    .io_mac_done    (uSystolicPE_244_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_244_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_244_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_244_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_244_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_244_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_244_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_0_5                     ), //i
    .io_ifm_dff     (ifm_dff_x_0_5                      ), //i
    .io_wght_sign   (wght_sign_x_5_0                    ), //i
    .io_randW       (randW_x_0_5[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_5_0[14:0]               ), //i
    .io_ofm         (ofm_x_5_1[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_244_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_244_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_244_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_244_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_244_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_244_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_244_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_244_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_244_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_244_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_244_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_244_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_244_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_245 (
    .io_mac_done    (uSystolicPE_245_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_245_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_245_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_245_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_245_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_245_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_245_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_0_6                     ), //i
    .io_ifm_dff     (ifm_dff_x_0_6                      ), //i
    .io_wght_sign   (wght_sign_x_6_0                    ), //i
    .io_randW       (randW_x_0_6[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_6_0[14:0]               ), //i
    .io_ofm         (ofm_x_6_1[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_245_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_245_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_245_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_245_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_245_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_245_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_245_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_245_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_245_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_245_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_245_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_245_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_245_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_246 (
    .io_mac_done    (uSystolicPE_246_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_246_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_246_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_246_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_246_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_246_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_246_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_0_7                     ), //i
    .io_ifm_dff     (ifm_dff_x_0_7                      ), //i
    .io_wght_sign   (wght_sign_x_7_0                    ), //i
    .io_randW       (randW_x_0_7[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_7_0[14:0]               ), //i
    .io_ofm         (ofm_x_7_1[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_246_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_246_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_246_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_246_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_246_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_246_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_246_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_246_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_246_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_246_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_246_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_246_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_246_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_247 (
    .io_mac_done    (uSystolicPE_247_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_247_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_247_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_247_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_247_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_247_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_247_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_0_8                     ), //i
    .io_ifm_dff     (ifm_dff_x_0_8                      ), //i
    .io_wght_sign   (wght_sign_x_8_0                    ), //i
    .io_randW       (randW_x_0_8[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_8_0[14:0]               ), //i
    .io_ofm         (ofm_x_8_1[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_247_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_247_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_247_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_247_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_247_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_247_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_247_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_247_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_247_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_247_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_247_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_247_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_247_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_248 (
    .io_mac_done    (uSystolicPE_248_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_248_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_248_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_248_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_248_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_248_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_248_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_0_9                     ), //i
    .io_ifm_dff     (ifm_dff_x_0_9                      ), //i
    .io_wght_sign   (wght_sign_x_9_0                    ), //i
    .io_randW       (randW_x_0_9[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_9_0[14:0]               ), //i
    .io_ofm         (ofm_x_9_1[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_248_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_248_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_248_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_248_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_248_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_248_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_248_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_248_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_248_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_248_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_248_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_248_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_248_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_249 (
    .io_mac_done    (uSystolicPE_249_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_249_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_249_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_249_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_249_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_249_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_249_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_0_10                    ), //i
    .io_ifm_dff     (ifm_dff_x_0_10                     ), //i
    .io_wght_sign   (wght_sign_x_10_0                   ), //i
    .io_randW       (randW_x_0_10[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_10_0[14:0]              ), //i
    .io_ofm         (ofm_x_10_1[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_249_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_249_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_249_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_249_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_249_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_249_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_249_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_249_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_249_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_249_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_249_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_249_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_249_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_250 (
    .io_mac_done    (uSystolicPE_250_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_250_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_250_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_250_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_250_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_250_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_250_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_0_11                    ), //i
    .io_ifm_dff     (ifm_dff_x_0_11                     ), //i
    .io_wght_sign   (wght_sign_x_11_0                   ), //i
    .io_randW       (randW_x_0_11[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_11_0[14:0]              ), //i
    .io_ofm         (ofm_x_11_1[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_250_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_250_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_250_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_250_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_250_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_250_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_250_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_250_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_250_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_250_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_250_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_250_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_250_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_251 (
    .io_mac_done    (uSystolicPE_251_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_251_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_251_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_251_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_251_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_251_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_251_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_0_12                    ), //i
    .io_ifm_dff     (ifm_dff_x_0_12                     ), //i
    .io_wght_sign   (wght_sign_x_12_0                   ), //i
    .io_randW       (randW_x_0_12[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_12_0[14:0]              ), //i
    .io_ofm         (ofm_x_12_1[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_251_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_251_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_251_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_251_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_251_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_251_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_251_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_251_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_251_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_251_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_251_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_251_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_251_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_252 (
    .io_mac_done    (uSystolicPE_252_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_252_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_252_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_252_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_252_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_252_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_252_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_0_13                    ), //i
    .io_ifm_dff     (ifm_dff_x_0_13                     ), //i
    .io_wght_sign   (wght_sign_x_13_0                   ), //i
    .io_randW       (randW_x_0_13[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_13_0[14:0]              ), //i
    .io_ofm         (ofm_x_13_1[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_252_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_252_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_252_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_252_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_252_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_252_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_252_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_252_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_252_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_252_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_252_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_252_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_252_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_253 (
    .io_mac_done    (uSystolicPE_253_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_253_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_253_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_253_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_253_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_253_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_253_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_0_14                    ), //i
    .io_ifm_dff     (ifm_dff_x_0_14                     ), //i
    .io_wght_sign   (wght_sign_x_14_0                   ), //i
    .io_randW       (randW_x_0_14[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_14_0[14:0]              ), //i
    .io_ofm         (ofm_x_14_1[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_253_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_253_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_253_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_253_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_253_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_253_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_253_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_253_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_253_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_253_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_253_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_253_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_253_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_254 (
    .io_mac_done    (uSystolicPE_254_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_254_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_254_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_254_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_254_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_254_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_254_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_0_15                    ), //i
    .io_ifm_dff     (ifm_dff_x_0_15                     ), //i
    .io_wght_sign   (wght_sign_x_15_0                   ), //i
    .io_randW       (randW_x_0_15[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_15_0[14:0]              ), //i
    .io_ofm         (ofm_x_15_1[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_254_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_254_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_254_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_254_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_254_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_254_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_254_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_254_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_254_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_254_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_254_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_254_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_254_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPEBorder uSystolicPEBorder_17 (
    .io_mac_done    (uSystolicPEBorder_17_io_mac_done        ), //i
    .io_enable_i    (uSystolicPEBorder_17_io_enable_i        ), //i
    .io_clear_i     (uSystolicPEBorder_17_io_clear_i         ), //i
    .io_enable_w    (uSystolicPEBorder_17_io_enable_w        ), //i
    .io_clear_w     (uSystolicPEBorder_17_io_clear_w         ), //i
    .io_enable_o    (uSystolicPEBorder_17_io_enable_o        ), //i
    .io_clear_o     (uSystolicPEBorder_17_io_clear_o         ), //i
    .io_ifm         (io_ifm_1[15:0]                          ), //i
    .io_wght_sign   (wght_sign_x_0_1                         ), //i
    .io_wght_abs    (wght_abs_x_0_1[14:0]                    ), //i
    .io_ofm         (ofm_x_0_2[31:0]                         ), //i
    .io_mac_done_d  (uSystolicPEBorder_17_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPEBorder_17_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPEBorder_17_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPEBorder_17_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPEBorder_17_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPEBorder_17_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPEBorder_17_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPEBorder_17_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPEBorder_17_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPEBorder_17_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPEBorder_17_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPEBorder_17_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPEBorder_17_io_ofm_d[31:0]     ), //o
    .clk            (clk                                     ), //i
    .reset          (reset                                   )  //i
  );
  uSystolicPE uSystolicPE_255 (
    .io_mac_done    (uSystolicPE_255_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_255_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_255_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_255_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_255_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_255_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_255_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_1_1                     ), //i
    .io_ifm_dff     (ifm_dff_x_1_1                      ), //i
    .io_wght_sign   (wght_sign_x_1_1                    ), //i
    .io_randW       (randW_x_1_1[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_1_1[14:0]               ), //i
    .io_ofm         (ofm_x_1_2[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_255_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_255_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_255_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_255_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_255_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_255_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_255_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_255_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_255_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_255_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_255_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_255_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_255_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_256 (
    .io_mac_done    (uSystolicPE_256_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_256_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_256_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_256_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_256_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_256_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_256_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_1_2                     ), //i
    .io_ifm_dff     (ifm_dff_x_1_2                      ), //i
    .io_wght_sign   (wght_sign_x_2_1                    ), //i
    .io_randW       (randW_x_1_2[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_2_1[14:0]               ), //i
    .io_ofm         (ofm_x_2_2[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_256_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_256_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_256_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_256_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_256_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_256_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_256_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_256_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_256_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_256_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_256_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_256_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_256_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_257 (
    .io_mac_done    (uSystolicPE_257_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_257_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_257_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_257_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_257_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_257_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_257_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_1_3                     ), //i
    .io_ifm_dff     (ifm_dff_x_1_3                      ), //i
    .io_wght_sign   (wght_sign_x_3_1                    ), //i
    .io_randW       (randW_x_1_3[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_3_1[14:0]               ), //i
    .io_ofm         (ofm_x_3_2[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_257_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_257_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_257_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_257_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_257_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_257_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_257_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_257_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_257_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_257_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_257_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_257_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_257_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_258 (
    .io_mac_done    (uSystolicPE_258_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_258_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_258_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_258_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_258_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_258_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_258_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_1_4                     ), //i
    .io_ifm_dff     (ifm_dff_x_1_4                      ), //i
    .io_wght_sign   (wght_sign_x_4_1                    ), //i
    .io_randW       (randW_x_1_4[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_4_1[14:0]               ), //i
    .io_ofm         (ofm_x_4_2[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_258_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_258_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_258_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_258_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_258_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_258_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_258_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_258_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_258_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_258_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_258_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_258_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_258_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_259 (
    .io_mac_done    (uSystolicPE_259_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_259_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_259_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_259_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_259_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_259_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_259_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_1_5                     ), //i
    .io_ifm_dff     (ifm_dff_x_1_5                      ), //i
    .io_wght_sign   (wght_sign_x_5_1                    ), //i
    .io_randW       (randW_x_1_5[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_5_1[14:0]               ), //i
    .io_ofm         (ofm_x_5_2[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_259_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_259_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_259_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_259_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_259_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_259_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_259_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_259_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_259_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_259_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_259_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_259_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_259_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_260 (
    .io_mac_done    (uSystolicPE_260_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_260_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_260_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_260_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_260_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_260_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_260_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_1_6                     ), //i
    .io_ifm_dff     (ifm_dff_x_1_6                      ), //i
    .io_wght_sign   (wght_sign_x_6_1                    ), //i
    .io_randW       (randW_x_1_6[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_6_1[14:0]               ), //i
    .io_ofm         (ofm_x_6_2[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_260_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_260_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_260_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_260_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_260_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_260_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_260_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_260_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_260_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_260_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_260_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_260_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_260_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_261 (
    .io_mac_done    (uSystolicPE_261_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_261_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_261_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_261_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_261_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_261_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_261_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_1_7                     ), //i
    .io_ifm_dff     (ifm_dff_x_1_7                      ), //i
    .io_wght_sign   (wght_sign_x_7_1                    ), //i
    .io_randW       (randW_x_1_7[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_7_1[14:0]               ), //i
    .io_ofm         (ofm_x_7_2[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_261_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_261_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_261_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_261_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_261_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_261_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_261_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_261_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_261_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_261_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_261_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_261_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_261_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_262 (
    .io_mac_done    (uSystolicPE_262_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_262_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_262_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_262_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_262_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_262_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_262_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_1_8                     ), //i
    .io_ifm_dff     (ifm_dff_x_1_8                      ), //i
    .io_wght_sign   (wght_sign_x_8_1                    ), //i
    .io_randW       (randW_x_1_8[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_8_1[14:0]               ), //i
    .io_ofm         (ofm_x_8_2[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_262_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_262_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_262_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_262_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_262_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_262_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_262_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_262_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_262_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_262_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_262_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_262_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_262_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_263 (
    .io_mac_done    (uSystolicPE_263_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_263_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_263_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_263_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_263_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_263_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_263_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_1_9                     ), //i
    .io_ifm_dff     (ifm_dff_x_1_9                      ), //i
    .io_wght_sign   (wght_sign_x_9_1                    ), //i
    .io_randW       (randW_x_1_9[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_9_1[14:0]               ), //i
    .io_ofm         (ofm_x_9_2[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_263_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_263_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_263_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_263_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_263_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_263_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_263_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_263_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_263_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_263_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_263_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_263_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_263_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_264 (
    .io_mac_done    (uSystolicPE_264_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_264_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_264_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_264_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_264_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_264_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_264_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_1_10                    ), //i
    .io_ifm_dff     (ifm_dff_x_1_10                     ), //i
    .io_wght_sign   (wght_sign_x_10_1                   ), //i
    .io_randW       (randW_x_1_10[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_10_1[14:0]              ), //i
    .io_ofm         (ofm_x_10_2[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_264_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_264_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_264_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_264_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_264_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_264_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_264_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_264_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_264_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_264_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_264_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_264_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_264_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_265 (
    .io_mac_done    (uSystolicPE_265_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_265_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_265_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_265_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_265_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_265_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_265_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_1_11                    ), //i
    .io_ifm_dff     (ifm_dff_x_1_11                     ), //i
    .io_wght_sign   (wght_sign_x_11_1                   ), //i
    .io_randW       (randW_x_1_11[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_11_1[14:0]              ), //i
    .io_ofm         (ofm_x_11_2[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_265_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_265_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_265_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_265_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_265_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_265_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_265_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_265_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_265_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_265_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_265_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_265_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_265_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_266 (
    .io_mac_done    (uSystolicPE_266_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_266_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_266_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_266_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_266_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_266_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_266_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_1_12                    ), //i
    .io_ifm_dff     (ifm_dff_x_1_12                     ), //i
    .io_wght_sign   (wght_sign_x_12_1                   ), //i
    .io_randW       (randW_x_1_12[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_12_1[14:0]              ), //i
    .io_ofm         (ofm_x_12_2[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_266_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_266_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_266_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_266_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_266_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_266_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_266_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_266_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_266_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_266_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_266_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_266_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_266_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_267 (
    .io_mac_done    (uSystolicPE_267_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_267_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_267_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_267_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_267_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_267_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_267_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_1_13                    ), //i
    .io_ifm_dff     (ifm_dff_x_1_13                     ), //i
    .io_wght_sign   (wght_sign_x_13_1                   ), //i
    .io_randW       (randW_x_1_13[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_13_1[14:0]              ), //i
    .io_ofm         (ofm_x_13_2[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_267_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_267_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_267_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_267_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_267_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_267_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_267_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_267_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_267_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_267_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_267_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_267_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_267_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_268 (
    .io_mac_done    (uSystolicPE_268_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_268_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_268_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_268_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_268_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_268_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_268_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_1_14                    ), //i
    .io_ifm_dff     (ifm_dff_x_1_14                     ), //i
    .io_wght_sign   (wght_sign_x_14_1                   ), //i
    .io_randW       (randW_x_1_14[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_14_1[14:0]              ), //i
    .io_ofm         (ofm_x_14_2[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_268_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_268_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_268_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_268_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_268_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_268_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_268_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_268_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_268_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_268_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_268_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_268_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_268_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_269 (
    .io_mac_done    (uSystolicPE_269_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_269_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_269_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_269_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_269_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_269_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_269_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_1_15                    ), //i
    .io_ifm_dff     (ifm_dff_x_1_15                     ), //i
    .io_wght_sign   (wght_sign_x_15_1                   ), //i
    .io_randW       (randW_x_1_15[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_15_1[14:0]              ), //i
    .io_ofm         (ofm_x_15_2[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_269_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_269_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_269_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_269_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_269_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_269_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_269_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_269_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_269_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_269_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_269_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_269_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_269_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPEBorder uSystolicPEBorder_18 (
    .io_mac_done    (uSystolicPEBorder_18_io_mac_done        ), //i
    .io_enable_i    (uSystolicPEBorder_18_io_enable_i        ), //i
    .io_clear_i     (uSystolicPEBorder_18_io_clear_i         ), //i
    .io_enable_w    (uSystolicPEBorder_18_io_enable_w        ), //i
    .io_clear_w     (uSystolicPEBorder_18_io_clear_w         ), //i
    .io_enable_o    (uSystolicPEBorder_18_io_enable_o        ), //i
    .io_clear_o     (uSystolicPEBorder_18_io_clear_o         ), //i
    .io_ifm         (io_ifm_2[15:0]                          ), //i
    .io_wght_sign   (wght_sign_x_0_2                         ), //i
    .io_wght_abs    (wght_abs_x_0_2[14:0]                    ), //i
    .io_ofm         (ofm_x_0_3[31:0]                         ), //i
    .io_mac_done_d  (uSystolicPEBorder_18_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPEBorder_18_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPEBorder_18_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPEBorder_18_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPEBorder_18_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPEBorder_18_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPEBorder_18_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPEBorder_18_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPEBorder_18_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPEBorder_18_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPEBorder_18_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPEBorder_18_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPEBorder_18_io_ofm_d[31:0]     ), //o
    .clk            (clk                                     ), //i
    .reset          (reset                                   )  //i
  );
  uSystolicPE uSystolicPE_270 (
    .io_mac_done    (uSystolicPE_270_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_270_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_270_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_270_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_270_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_270_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_270_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_2_1                     ), //i
    .io_ifm_dff     (ifm_dff_x_2_1                      ), //i
    .io_wght_sign   (wght_sign_x_1_2                    ), //i
    .io_randW       (randW_x_2_1[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_1_2[14:0]               ), //i
    .io_ofm         (ofm_x_1_3[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_270_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_270_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_270_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_270_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_270_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_270_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_270_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_270_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_270_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_270_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_270_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_270_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_270_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_271 (
    .io_mac_done    (uSystolicPE_271_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_271_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_271_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_271_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_271_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_271_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_271_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_2_2                     ), //i
    .io_ifm_dff     (ifm_dff_x_2_2                      ), //i
    .io_wght_sign   (wght_sign_x_2_2                    ), //i
    .io_randW       (randW_x_2_2[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_2_2[14:0]               ), //i
    .io_ofm         (ofm_x_2_3[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_271_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_271_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_271_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_271_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_271_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_271_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_271_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_271_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_271_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_271_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_271_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_271_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_271_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_272 (
    .io_mac_done    (uSystolicPE_272_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_272_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_272_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_272_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_272_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_272_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_272_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_2_3                     ), //i
    .io_ifm_dff     (ifm_dff_x_2_3                      ), //i
    .io_wght_sign   (wght_sign_x_3_2                    ), //i
    .io_randW       (randW_x_2_3[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_3_2[14:0]               ), //i
    .io_ofm         (ofm_x_3_3[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_272_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_272_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_272_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_272_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_272_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_272_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_272_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_272_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_272_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_272_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_272_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_272_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_272_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_273 (
    .io_mac_done    (uSystolicPE_273_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_273_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_273_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_273_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_273_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_273_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_273_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_2_4                     ), //i
    .io_ifm_dff     (ifm_dff_x_2_4                      ), //i
    .io_wght_sign   (wght_sign_x_4_2                    ), //i
    .io_randW       (randW_x_2_4[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_4_2[14:0]               ), //i
    .io_ofm         (ofm_x_4_3[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_273_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_273_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_273_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_273_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_273_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_273_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_273_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_273_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_273_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_273_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_273_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_273_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_273_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_274 (
    .io_mac_done    (uSystolicPE_274_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_274_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_274_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_274_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_274_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_274_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_274_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_2_5                     ), //i
    .io_ifm_dff     (ifm_dff_x_2_5                      ), //i
    .io_wght_sign   (wght_sign_x_5_2                    ), //i
    .io_randW       (randW_x_2_5[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_5_2[14:0]               ), //i
    .io_ofm         (ofm_x_5_3[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_274_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_274_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_274_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_274_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_274_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_274_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_274_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_274_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_274_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_274_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_274_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_274_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_274_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_275 (
    .io_mac_done    (uSystolicPE_275_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_275_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_275_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_275_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_275_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_275_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_275_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_2_6                     ), //i
    .io_ifm_dff     (ifm_dff_x_2_6                      ), //i
    .io_wght_sign   (wght_sign_x_6_2                    ), //i
    .io_randW       (randW_x_2_6[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_6_2[14:0]               ), //i
    .io_ofm         (ofm_x_6_3[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_275_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_275_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_275_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_275_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_275_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_275_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_275_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_275_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_275_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_275_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_275_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_275_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_275_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_276 (
    .io_mac_done    (uSystolicPE_276_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_276_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_276_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_276_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_276_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_276_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_276_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_2_7                     ), //i
    .io_ifm_dff     (ifm_dff_x_2_7                      ), //i
    .io_wght_sign   (wght_sign_x_7_2                    ), //i
    .io_randW       (randW_x_2_7[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_7_2[14:0]               ), //i
    .io_ofm         (ofm_x_7_3[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_276_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_276_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_276_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_276_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_276_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_276_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_276_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_276_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_276_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_276_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_276_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_276_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_276_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_277 (
    .io_mac_done    (uSystolicPE_277_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_277_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_277_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_277_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_277_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_277_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_277_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_2_8                     ), //i
    .io_ifm_dff     (ifm_dff_x_2_8                      ), //i
    .io_wght_sign   (wght_sign_x_8_2                    ), //i
    .io_randW       (randW_x_2_8[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_8_2[14:0]               ), //i
    .io_ofm         (ofm_x_8_3[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_277_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_277_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_277_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_277_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_277_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_277_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_277_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_277_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_277_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_277_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_277_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_277_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_277_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_278 (
    .io_mac_done    (uSystolicPE_278_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_278_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_278_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_278_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_278_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_278_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_278_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_2_9                     ), //i
    .io_ifm_dff     (ifm_dff_x_2_9                      ), //i
    .io_wght_sign   (wght_sign_x_9_2                    ), //i
    .io_randW       (randW_x_2_9[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_9_2[14:0]               ), //i
    .io_ofm         (ofm_x_9_3[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_278_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_278_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_278_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_278_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_278_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_278_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_278_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_278_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_278_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_278_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_278_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_278_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_278_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_279 (
    .io_mac_done    (uSystolicPE_279_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_279_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_279_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_279_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_279_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_279_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_279_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_2_10                    ), //i
    .io_ifm_dff     (ifm_dff_x_2_10                     ), //i
    .io_wght_sign   (wght_sign_x_10_2                   ), //i
    .io_randW       (randW_x_2_10[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_10_2[14:0]              ), //i
    .io_ofm         (ofm_x_10_3[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_279_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_279_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_279_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_279_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_279_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_279_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_279_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_279_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_279_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_279_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_279_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_279_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_279_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_280 (
    .io_mac_done    (uSystolicPE_280_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_280_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_280_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_280_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_280_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_280_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_280_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_2_11                    ), //i
    .io_ifm_dff     (ifm_dff_x_2_11                     ), //i
    .io_wght_sign   (wght_sign_x_11_2                   ), //i
    .io_randW       (randW_x_2_11[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_11_2[14:0]              ), //i
    .io_ofm         (ofm_x_11_3[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_280_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_280_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_280_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_280_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_280_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_280_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_280_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_280_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_280_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_280_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_280_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_280_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_280_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_281 (
    .io_mac_done    (uSystolicPE_281_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_281_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_281_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_281_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_281_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_281_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_281_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_2_12                    ), //i
    .io_ifm_dff     (ifm_dff_x_2_12                     ), //i
    .io_wght_sign   (wght_sign_x_12_2                   ), //i
    .io_randW       (randW_x_2_12[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_12_2[14:0]              ), //i
    .io_ofm         (ofm_x_12_3[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_281_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_281_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_281_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_281_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_281_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_281_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_281_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_281_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_281_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_281_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_281_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_281_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_281_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_282 (
    .io_mac_done    (uSystolicPE_282_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_282_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_282_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_282_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_282_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_282_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_282_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_2_13                    ), //i
    .io_ifm_dff     (ifm_dff_x_2_13                     ), //i
    .io_wght_sign   (wght_sign_x_13_2                   ), //i
    .io_randW       (randW_x_2_13[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_13_2[14:0]              ), //i
    .io_ofm         (ofm_x_13_3[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_282_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_282_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_282_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_282_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_282_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_282_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_282_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_282_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_282_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_282_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_282_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_282_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_282_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_283 (
    .io_mac_done    (uSystolicPE_283_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_283_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_283_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_283_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_283_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_283_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_283_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_2_14                    ), //i
    .io_ifm_dff     (ifm_dff_x_2_14                     ), //i
    .io_wght_sign   (wght_sign_x_14_2                   ), //i
    .io_randW       (randW_x_2_14[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_14_2[14:0]              ), //i
    .io_ofm         (ofm_x_14_3[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_283_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_283_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_283_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_283_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_283_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_283_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_283_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_283_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_283_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_283_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_283_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_283_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_283_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_284 (
    .io_mac_done    (uSystolicPE_284_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_284_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_284_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_284_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_284_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_284_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_284_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_2_15                    ), //i
    .io_ifm_dff     (ifm_dff_x_2_15                     ), //i
    .io_wght_sign   (wght_sign_x_15_2                   ), //i
    .io_randW       (randW_x_2_15[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_15_2[14:0]              ), //i
    .io_ofm         (ofm_x_15_3[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_284_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_284_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_284_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_284_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_284_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_284_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_284_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_284_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_284_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_284_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_284_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_284_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_284_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPEBorder uSystolicPEBorder_19 (
    .io_mac_done    (uSystolicPEBorder_19_io_mac_done        ), //i
    .io_enable_i    (uSystolicPEBorder_19_io_enable_i        ), //i
    .io_clear_i     (uSystolicPEBorder_19_io_clear_i         ), //i
    .io_enable_w    (uSystolicPEBorder_19_io_enable_w        ), //i
    .io_clear_w     (uSystolicPEBorder_19_io_clear_w         ), //i
    .io_enable_o    (uSystolicPEBorder_19_io_enable_o        ), //i
    .io_clear_o     (uSystolicPEBorder_19_io_clear_o         ), //i
    .io_ifm         (io_ifm_3[15:0]                          ), //i
    .io_wght_sign   (wght_sign_x_0_3                         ), //i
    .io_wght_abs    (wght_abs_x_0_3[14:0]                    ), //i
    .io_ofm         (ofm_x_0_4[31:0]                         ), //i
    .io_mac_done_d  (uSystolicPEBorder_19_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPEBorder_19_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPEBorder_19_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPEBorder_19_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPEBorder_19_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPEBorder_19_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPEBorder_19_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPEBorder_19_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPEBorder_19_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPEBorder_19_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPEBorder_19_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPEBorder_19_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPEBorder_19_io_ofm_d[31:0]     ), //o
    .clk            (clk                                     ), //i
    .reset          (reset                                   )  //i
  );
  uSystolicPE uSystolicPE_285 (
    .io_mac_done    (uSystolicPE_285_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_285_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_285_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_285_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_285_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_285_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_285_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_3_1                     ), //i
    .io_ifm_dff     (ifm_dff_x_3_1                      ), //i
    .io_wght_sign   (wght_sign_x_1_3                    ), //i
    .io_randW       (randW_x_3_1[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_1_3[14:0]               ), //i
    .io_ofm         (ofm_x_1_4[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_285_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_285_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_285_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_285_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_285_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_285_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_285_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_285_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_285_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_285_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_285_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_285_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_285_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_286 (
    .io_mac_done    (uSystolicPE_286_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_286_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_286_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_286_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_286_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_286_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_286_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_3_2                     ), //i
    .io_ifm_dff     (ifm_dff_x_3_2                      ), //i
    .io_wght_sign   (wght_sign_x_2_3                    ), //i
    .io_randW       (randW_x_3_2[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_2_3[14:0]               ), //i
    .io_ofm         (ofm_x_2_4[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_286_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_286_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_286_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_286_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_286_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_286_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_286_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_286_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_286_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_286_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_286_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_286_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_286_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_287 (
    .io_mac_done    (uSystolicPE_287_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_287_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_287_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_287_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_287_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_287_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_287_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_3_3                     ), //i
    .io_ifm_dff     (ifm_dff_x_3_3                      ), //i
    .io_wght_sign   (wght_sign_x_3_3                    ), //i
    .io_randW       (randW_x_3_3[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_3_3[14:0]               ), //i
    .io_ofm         (ofm_x_3_4[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_287_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_287_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_287_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_287_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_287_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_287_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_287_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_287_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_287_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_287_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_287_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_287_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_287_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_288 (
    .io_mac_done    (uSystolicPE_288_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_288_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_288_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_288_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_288_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_288_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_288_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_3_4                     ), //i
    .io_ifm_dff     (ifm_dff_x_3_4                      ), //i
    .io_wght_sign   (wght_sign_x_4_3                    ), //i
    .io_randW       (randW_x_3_4[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_4_3[14:0]               ), //i
    .io_ofm         (ofm_x_4_4[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_288_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_288_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_288_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_288_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_288_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_288_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_288_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_288_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_288_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_288_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_288_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_288_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_288_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_289 (
    .io_mac_done    (uSystolicPE_289_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_289_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_289_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_289_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_289_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_289_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_289_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_3_5                     ), //i
    .io_ifm_dff     (ifm_dff_x_3_5                      ), //i
    .io_wght_sign   (wght_sign_x_5_3                    ), //i
    .io_randW       (randW_x_3_5[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_5_3[14:0]               ), //i
    .io_ofm         (ofm_x_5_4[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_289_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_289_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_289_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_289_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_289_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_289_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_289_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_289_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_289_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_289_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_289_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_289_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_289_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_290 (
    .io_mac_done    (uSystolicPE_290_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_290_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_290_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_290_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_290_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_290_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_290_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_3_6                     ), //i
    .io_ifm_dff     (ifm_dff_x_3_6                      ), //i
    .io_wght_sign   (wght_sign_x_6_3                    ), //i
    .io_randW       (randW_x_3_6[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_6_3[14:0]               ), //i
    .io_ofm         (ofm_x_6_4[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_290_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_290_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_290_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_290_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_290_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_290_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_290_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_290_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_290_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_290_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_290_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_290_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_290_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_291 (
    .io_mac_done    (uSystolicPE_291_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_291_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_291_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_291_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_291_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_291_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_291_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_3_7                     ), //i
    .io_ifm_dff     (ifm_dff_x_3_7                      ), //i
    .io_wght_sign   (wght_sign_x_7_3                    ), //i
    .io_randW       (randW_x_3_7[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_7_3[14:0]               ), //i
    .io_ofm         (ofm_x_7_4[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_291_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_291_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_291_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_291_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_291_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_291_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_291_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_291_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_291_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_291_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_291_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_291_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_291_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_292 (
    .io_mac_done    (uSystolicPE_292_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_292_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_292_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_292_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_292_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_292_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_292_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_3_8                     ), //i
    .io_ifm_dff     (ifm_dff_x_3_8                      ), //i
    .io_wght_sign   (wght_sign_x_8_3                    ), //i
    .io_randW       (randW_x_3_8[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_8_3[14:0]               ), //i
    .io_ofm         (ofm_x_8_4[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_292_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_292_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_292_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_292_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_292_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_292_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_292_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_292_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_292_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_292_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_292_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_292_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_292_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_293 (
    .io_mac_done    (uSystolicPE_293_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_293_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_293_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_293_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_293_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_293_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_293_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_3_9                     ), //i
    .io_ifm_dff     (ifm_dff_x_3_9                      ), //i
    .io_wght_sign   (wght_sign_x_9_3                    ), //i
    .io_randW       (randW_x_3_9[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_9_3[14:0]               ), //i
    .io_ofm         (ofm_x_9_4[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_293_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_293_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_293_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_293_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_293_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_293_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_293_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_293_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_293_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_293_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_293_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_293_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_293_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_294 (
    .io_mac_done    (uSystolicPE_294_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_294_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_294_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_294_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_294_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_294_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_294_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_3_10                    ), //i
    .io_ifm_dff     (ifm_dff_x_3_10                     ), //i
    .io_wght_sign   (wght_sign_x_10_3                   ), //i
    .io_randW       (randW_x_3_10[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_10_3[14:0]              ), //i
    .io_ofm         (ofm_x_10_4[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_294_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_294_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_294_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_294_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_294_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_294_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_294_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_294_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_294_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_294_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_294_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_294_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_294_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_295 (
    .io_mac_done    (uSystolicPE_295_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_295_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_295_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_295_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_295_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_295_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_295_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_3_11                    ), //i
    .io_ifm_dff     (ifm_dff_x_3_11                     ), //i
    .io_wght_sign   (wght_sign_x_11_3                   ), //i
    .io_randW       (randW_x_3_11[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_11_3[14:0]              ), //i
    .io_ofm         (ofm_x_11_4[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_295_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_295_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_295_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_295_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_295_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_295_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_295_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_295_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_295_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_295_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_295_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_295_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_295_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_296 (
    .io_mac_done    (uSystolicPE_296_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_296_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_296_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_296_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_296_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_296_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_296_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_3_12                    ), //i
    .io_ifm_dff     (ifm_dff_x_3_12                     ), //i
    .io_wght_sign   (wght_sign_x_12_3                   ), //i
    .io_randW       (randW_x_3_12[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_12_3[14:0]              ), //i
    .io_ofm         (ofm_x_12_4[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_296_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_296_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_296_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_296_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_296_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_296_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_296_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_296_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_296_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_296_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_296_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_296_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_296_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_297 (
    .io_mac_done    (uSystolicPE_297_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_297_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_297_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_297_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_297_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_297_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_297_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_3_13                    ), //i
    .io_ifm_dff     (ifm_dff_x_3_13                     ), //i
    .io_wght_sign   (wght_sign_x_13_3                   ), //i
    .io_randW       (randW_x_3_13[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_13_3[14:0]              ), //i
    .io_ofm         (ofm_x_13_4[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_297_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_297_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_297_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_297_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_297_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_297_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_297_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_297_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_297_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_297_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_297_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_297_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_297_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_298 (
    .io_mac_done    (uSystolicPE_298_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_298_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_298_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_298_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_298_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_298_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_298_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_3_14                    ), //i
    .io_ifm_dff     (ifm_dff_x_3_14                     ), //i
    .io_wght_sign   (wght_sign_x_14_3                   ), //i
    .io_randW       (randW_x_3_14[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_14_3[14:0]              ), //i
    .io_ofm         (ofm_x_14_4[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_298_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_298_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_298_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_298_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_298_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_298_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_298_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_298_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_298_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_298_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_298_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_298_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_298_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_299 (
    .io_mac_done    (uSystolicPE_299_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_299_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_299_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_299_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_299_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_299_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_299_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_3_15                    ), //i
    .io_ifm_dff     (ifm_dff_x_3_15                     ), //i
    .io_wght_sign   (wght_sign_x_15_3                   ), //i
    .io_randW       (randW_x_3_15[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_15_3[14:0]              ), //i
    .io_ofm         (ofm_x_15_4[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_299_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_299_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_299_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_299_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_299_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_299_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_299_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_299_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_299_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_299_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_299_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_299_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_299_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPEBorder uSystolicPEBorder_20 (
    .io_mac_done    (uSystolicPEBorder_20_io_mac_done        ), //i
    .io_enable_i    (uSystolicPEBorder_20_io_enable_i        ), //i
    .io_clear_i     (uSystolicPEBorder_20_io_clear_i         ), //i
    .io_enable_w    (uSystolicPEBorder_20_io_enable_w        ), //i
    .io_clear_w     (uSystolicPEBorder_20_io_clear_w         ), //i
    .io_enable_o    (uSystolicPEBorder_20_io_enable_o        ), //i
    .io_clear_o     (uSystolicPEBorder_20_io_clear_o         ), //i
    .io_ifm         (io_ifm_4[15:0]                          ), //i
    .io_wght_sign   (wght_sign_x_0_4                         ), //i
    .io_wght_abs    (wght_abs_x_0_4[14:0]                    ), //i
    .io_ofm         (ofm_x_0_5[31:0]                         ), //i
    .io_mac_done_d  (uSystolicPEBorder_20_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPEBorder_20_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPEBorder_20_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPEBorder_20_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPEBorder_20_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPEBorder_20_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPEBorder_20_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPEBorder_20_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPEBorder_20_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPEBorder_20_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPEBorder_20_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPEBorder_20_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPEBorder_20_io_ofm_d[31:0]     ), //o
    .clk            (clk                                     ), //i
    .reset          (reset                                   )  //i
  );
  uSystolicPE uSystolicPE_300 (
    .io_mac_done    (uSystolicPE_300_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_300_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_300_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_300_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_300_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_300_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_300_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_4_1                     ), //i
    .io_ifm_dff     (ifm_dff_x_4_1                      ), //i
    .io_wght_sign   (wght_sign_x_1_4                    ), //i
    .io_randW       (randW_x_4_1[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_1_4[14:0]               ), //i
    .io_ofm         (ofm_x_1_5[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_300_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_300_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_300_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_300_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_300_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_300_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_300_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_300_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_300_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_300_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_300_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_300_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_300_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_301 (
    .io_mac_done    (uSystolicPE_301_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_301_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_301_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_301_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_301_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_301_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_301_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_4_2                     ), //i
    .io_ifm_dff     (ifm_dff_x_4_2                      ), //i
    .io_wght_sign   (wght_sign_x_2_4                    ), //i
    .io_randW       (randW_x_4_2[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_2_4[14:0]               ), //i
    .io_ofm         (ofm_x_2_5[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_301_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_301_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_301_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_301_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_301_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_301_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_301_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_301_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_301_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_301_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_301_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_301_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_301_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_302 (
    .io_mac_done    (uSystolicPE_302_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_302_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_302_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_302_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_302_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_302_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_302_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_4_3                     ), //i
    .io_ifm_dff     (ifm_dff_x_4_3                      ), //i
    .io_wght_sign   (wght_sign_x_3_4                    ), //i
    .io_randW       (randW_x_4_3[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_3_4[14:0]               ), //i
    .io_ofm         (ofm_x_3_5[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_302_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_302_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_302_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_302_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_302_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_302_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_302_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_302_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_302_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_302_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_302_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_302_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_302_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_303 (
    .io_mac_done    (uSystolicPE_303_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_303_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_303_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_303_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_303_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_303_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_303_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_4_4                     ), //i
    .io_ifm_dff     (ifm_dff_x_4_4                      ), //i
    .io_wght_sign   (wght_sign_x_4_4                    ), //i
    .io_randW       (randW_x_4_4[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_4_4[14:0]               ), //i
    .io_ofm         (ofm_x_4_5[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_303_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_303_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_303_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_303_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_303_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_303_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_303_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_303_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_303_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_303_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_303_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_303_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_303_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_304 (
    .io_mac_done    (uSystolicPE_304_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_304_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_304_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_304_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_304_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_304_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_304_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_4_5                     ), //i
    .io_ifm_dff     (ifm_dff_x_4_5                      ), //i
    .io_wght_sign   (wght_sign_x_5_4                    ), //i
    .io_randW       (randW_x_4_5[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_5_4[14:0]               ), //i
    .io_ofm         (ofm_x_5_5[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_304_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_304_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_304_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_304_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_304_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_304_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_304_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_304_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_304_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_304_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_304_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_304_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_304_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_305 (
    .io_mac_done    (uSystolicPE_305_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_305_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_305_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_305_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_305_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_305_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_305_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_4_6                     ), //i
    .io_ifm_dff     (ifm_dff_x_4_6                      ), //i
    .io_wght_sign   (wght_sign_x_6_4                    ), //i
    .io_randW       (randW_x_4_6[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_6_4[14:0]               ), //i
    .io_ofm         (ofm_x_6_5[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_305_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_305_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_305_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_305_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_305_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_305_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_305_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_305_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_305_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_305_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_305_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_305_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_305_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_306 (
    .io_mac_done    (uSystolicPE_306_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_306_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_306_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_306_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_306_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_306_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_306_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_4_7                     ), //i
    .io_ifm_dff     (ifm_dff_x_4_7                      ), //i
    .io_wght_sign   (wght_sign_x_7_4                    ), //i
    .io_randW       (randW_x_4_7[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_7_4[14:0]               ), //i
    .io_ofm         (ofm_x_7_5[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_306_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_306_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_306_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_306_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_306_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_306_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_306_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_306_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_306_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_306_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_306_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_306_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_306_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_307 (
    .io_mac_done    (uSystolicPE_307_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_307_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_307_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_307_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_307_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_307_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_307_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_4_8                     ), //i
    .io_ifm_dff     (ifm_dff_x_4_8                      ), //i
    .io_wght_sign   (wght_sign_x_8_4                    ), //i
    .io_randW       (randW_x_4_8[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_8_4[14:0]               ), //i
    .io_ofm         (ofm_x_8_5[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_307_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_307_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_307_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_307_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_307_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_307_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_307_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_307_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_307_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_307_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_307_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_307_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_307_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_308 (
    .io_mac_done    (uSystolicPE_308_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_308_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_308_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_308_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_308_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_308_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_308_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_4_9                     ), //i
    .io_ifm_dff     (ifm_dff_x_4_9                      ), //i
    .io_wght_sign   (wght_sign_x_9_4                    ), //i
    .io_randW       (randW_x_4_9[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_9_4[14:0]               ), //i
    .io_ofm         (ofm_x_9_5[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_308_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_308_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_308_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_308_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_308_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_308_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_308_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_308_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_308_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_308_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_308_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_308_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_308_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_309 (
    .io_mac_done    (uSystolicPE_309_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_309_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_309_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_309_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_309_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_309_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_309_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_4_10                    ), //i
    .io_ifm_dff     (ifm_dff_x_4_10                     ), //i
    .io_wght_sign   (wght_sign_x_10_4                   ), //i
    .io_randW       (randW_x_4_10[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_10_4[14:0]              ), //i
    .io_ofm         (ofm_x_10_5[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_309_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_309_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_309_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_309_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_309_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_309_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_309_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_309_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_309_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_309_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_309_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_309_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_309_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_310 (
    .io_mac_done    (uSystolicPE_310_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_310_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_310_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_310_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_310_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_310_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_310_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_4_11                    ), //i
    .io_ifm_dff     (ifm_dff_x_4_11                     ), //i
    .io_wght_sign   (wght_sign_x_11_4                   ), //i
    .io_randW       (randW_x_4_11[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_11_4[14:0]              ), //i
    .io_ofm         (ofm_x_11_5[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_310_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_310_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_310_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_310_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_310_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_310_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_310_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_310_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_310_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_310_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_310_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_310_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_310_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_311 (
    .io_mac_done    (uSystolicPE_311_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_311_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_311_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_311_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_311_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_311_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_311_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_4_12                    ), //i
    .io_ifm_dff     (ifm_dff_x_4_12                     ), //i
    .io_wght_sign   (wght_sign_x_12_4                   ), //i
    .io_randW       (randW_x_4_12[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_12_4[14:0]              ), //i
    .io_ofm         (ofm_x_12_5[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_311_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_311_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_311_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_311_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_311_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_311_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_311_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_311_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_311_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_311_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_311_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_311_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_311_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_312 (
    .io_mac_done    (uSystolicPE_312_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_312_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_312_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_312_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_312_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_312_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_312_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_4_13                    ), //i
    .io_ifm_dff     (ifm_dff_x_4_13                     ), //i
    .io_wght_sign   (wght_sign_x_13_4                   ), //i
    .io_randW       (randW_x_4_13[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_13_4[14:0]              ), //i
    .io_ofm         (ofm_x_13_5[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_312_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_312_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_312_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_312_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_312_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_312_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_312_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_312_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_312_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_312_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_312_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_312_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_312_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_313 (
    .io_mac_done    (uSystolicPE_313_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_313_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_313_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_313_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_313_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_313_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_313_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_4_14                    ), //i
    .io_ifm_dff     (ifm_dff_x_4_14                     ), //i
    .io_wght_sign   (wght_sign_x_14_4                   ), //i
    .io_randW       (randW_x_4_14[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_14_4[14:0]              ), //i
    .io_ofm         (ofm_x_14_5[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_313_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_313_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_313_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_313_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_313_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_313_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_313_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_313_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_313_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_313_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_313_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_313_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_313_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_314 (
    .io_mac_done    (uSystolicPE_314_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_314_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_314_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_314_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_314_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_314_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_314_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_4_15                    ), //i
    .io_ifm_dff     (ifm_dff_x_4_15                     ), //i
    .io_wght_sign   (wght_sign_x_15_4                   ), //i
    .io_randW       (randW_x_4_15[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_15_4[14:0]              ), //i
    .io_ofm         (ofm_x_15_5[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_314_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_314_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_314_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_314_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_314_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_314_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_314_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_314_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_314_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_314_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_314_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_314_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_314_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPEBorder uSystolicPEBorder_21 (
    .io_mac_done    (uSystolicPEBorder_21_io_mac_done        ), //i
    .io_enable_i    (uSystolicPEBorder_21_io_enable_i        ), //i
    .io_clear_i     (uSystolicPEBorder_21_io_clear_i         ), //i
    .io_enable_w    (uSystolicPEBorder_21_io_enable_w        ), //i
    .io_clear_w     (uSystolicPEBorder_21_io_clear_w         ), //i
    .io_enable_o    (uSystolicPEBorder_21_io_enable_o        ), //i
    .io_clear_o     (uSystolicPEBorder_21_io_clear_o         ), //i
    .io_ifm         (io_ifm_5[15:0]                          ), //i
    .io_wght_sign   (wght_sign_x_0_5                         ), //i
    .io_wght_abs    (wght_abs_x_0_5[14:0]                    ), //i
    .io_ofm         (ofm_x_0_6[31:0]                         ), //i
    .io_mac_done_d  (uSystolicPEBorder_21_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPEBorder_21_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPEBorder_21_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPEBorder_21_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPEBorder_21_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPEBorder_21_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPEBorder_21_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPEBorder_21_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPEBorder_21_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPEBorder_21_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPEBorder_21_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPEBorder_21_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPEBorder_21_io_ofm_d[31:0]     ), //o
    .clk            (clk                                     ), //i
    .reset          (reset                                   )  //i
  );
  uSystolicPE uSystolicPE_315 (
    .io_mac_done    (uSystolicPE_315_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_315_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_315_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_315_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_315_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_315_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_315_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_5_1                     ), //i
    .io_ifm_dff     (ifm_dff_x_5_1                      ), //i
    .io_wght_sign   (wght_sign_x_1_5                    ), //i
    .io_randW       (randW_x_5_1[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_1_5[14:0]               ), //i
    .io_ofm         (ofm_x_1_6[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_315_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_315_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_315_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_315_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_315_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_315_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_315_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_315_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_315_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_315_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_315_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_315_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_315_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_316 (
    .io_mac_done    (uSystolicPE_316_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_316_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_316_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_316_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_316_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_316_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_316_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_5_2                     ), //i
    .io_ifm_dff     (ifm_dff_x_5_2                      ), //i
    .io_wght_sign   (wght_sign_x_2_5                    ), //i
    .io_randW       (randW_x_5_2[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_2_5[14:0]               ), //i
    .io_ofm         (ofm_x_2_6[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_316_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_316_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_316_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_316_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_316_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_316_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_316_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_316_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_316_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_316_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_316_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_316_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_316_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_317 (
    .io_mac_done    (uSystolicPE_317_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_317_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_317_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_317_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_317_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_317_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_317_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_5_3                     ), //i
    .io_ifm_dff     (ifm_dff_x_5_3                      ), //i
    .io_wght_sign   (wght_sign_x_3_5                    ), //i
    .io_randW       (randW_x_5_3[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_3_5[14:0]               ), //i
    .io_ofm         (ofm_x_3_6[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_317_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_317_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_317_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_317_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_317_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_317_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_317_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_317_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_317_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_317_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_317_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_317_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_317_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_318 (
    .io_mac_done    (uSystolicPE_318_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_318_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_318_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_318_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_318_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_318_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_318_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_5_4                     ), //i
    .io_ifm_dff     (ifm_dff_x_5_4                      ), //i
    .io_wght_sign   (wght_sign_x_4_5                    ), //i
    .io_randW       (randW_x_5_4[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_4_5[14:0]               ), //i
    .io_ofm         (ofm_x_4_6[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_318_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_318_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_318_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_318_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_318_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_318_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_318_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_318_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_318_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_318_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_318_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_318_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_318_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_319 (
    .io_mac_done    (uSystolicPE_319_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_319_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_319_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_319_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_319_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_319_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_319_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_5_5                     ), //i
    .io_ifm_dff     (ifm_dff_x_5_5                      ), //i
    .io_wght_sign   (wght_sign_x_5_5                    ), //i
    .io_randW       (randW_x_5_5[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_5_5[14:0]               ), //i
    .io_ofm         (ofm_x_5_6[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_319_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_319_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_319_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_319_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_319_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_319_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_319_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_319_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_319_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_319_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_319_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_319_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_319_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_320 (
    .io_mac_done    (uSystolicPE_320_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_320_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_320_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_320_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_320_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_320_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_320_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_5_6                     ), //i
    .io_ifm_dff     (ifm_dff_x_5_6                      ), //i
    .io_wght_sign   (wght_sign_x_6_5                    ), //i
    .io_randW       (randW_x_5_6[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_6_5[14:0]               ), //i
    .io_ofm         (ofm_x_6_6[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_320_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_320_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_320_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_320_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_320_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_320_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_320_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_320_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_320_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_320_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_320_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_320_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_320_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_321 (
    .io_mac_done    (uSystolicPE_321_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_321_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_321_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_321_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_321_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_321_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_321_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_5_7                     ), //i
    .io_ifm_dff     (ifm_dff_x_5_7                      ), //i
    .io_wght_sign   (wght_sign_x_7_5                    ), //i
    .io_randW       (randW_x_5_7[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_7_5[14:0]               ), //i
    .io_ofm         (ofm_x_7_6[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_321_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_321_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_321_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_321_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_321_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_321_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_321_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_321_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_321_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_321_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_321_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_321_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_321_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_322 (
    .io_mac_done    (uSystolicPE_322_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_322_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_322_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_322_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_322_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_322_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_322_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_5_8                     ), //i
    .io_ifm_dff     (ifm_dff_x_5_8                      ), //i
    .io_wght_sign   (wght_sign_x_8_5                    ), //i
    .io_randW       (randW_x_5_8[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_8_5[14:0]               ), //i
    .io_ofm         (ofm_x_8_6[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_322_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_322_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_322_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_322_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_322_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_322_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_322_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_322_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_322_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_322_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_322_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_322_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_322_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_323 (
    .io_mac_done    (uSystolicPE_323_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_323_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_323_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_323_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_323_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_323_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_323_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_5_9                     ), //i
    .io_ifm_dff     (ifm_dff_x_5_9                      ), //i
    .io_wght_sign   (wght_sign_x_9_5                    ), //i
    .io_randW       (randW_x_5_9[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_9_5[14:0]               ), //i
    .io_ofm         (ofm_x_9_6[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_323_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_323_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_323_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_323_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_323_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_323_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_323_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_323_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_323_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_323_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_323_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_323_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_323_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_324 (
    .io_mac_done    (uSystolicPE_324_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_324_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_324_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_324_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_324_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_324_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_324_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_5_10                    ), //i
    .io_ifm_dff     (ifm_dff_x_5_10                     ), //i
    .io_wght_sign   (wght_sign_x_10_5                   ), //i
    .io_randW       (randW_x_5_10[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_10_5[14:0]              ), //i
    .io_ofm         (ofm_x_10_6[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_324_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_324_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_324_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_324_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_324_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_324_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_324_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_324_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_324_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_324_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_324_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_324_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_324_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_325 (
    .io_mac_done    (uSystolicPE_325_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_325_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_325_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_325_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_325_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_325_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_325_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_5_11                    ), //i
    .io_ifm_dff     (ifm_dff_x_5_11                     ), //i
    .io_wght_sign   (wght_sign_x_11_5                   ), //i
    .io_randW       (randW_x_5_11[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_11_5[14:0]              ), //i
    .io_ofm         (ofm_x_11_6[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_325_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_325_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_325_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_325_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_325_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_325_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_325_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_325_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_325_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_325_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_325_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_325_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_325_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_326 (
    .io_mac_done    (uSystolicPE_326_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_326_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_326_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_326_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_326_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_326_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_326_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_5_12                    ), //i
    .io_ifm_dff     (ifm_dff_x_5_12                     ), //i
    .io_wght_sign   (wght_sign_x_12_5                   ), //i
    .io_randW       (randW_x_5_12[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_12_5[14:0]              ), //i
    .io_ofm         (ofm_x_12_6[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_326_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_326_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_326_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_326_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_326_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_326_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_326_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_326_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_326_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_326_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_326_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_326_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_326_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_327 (
    .io_mac_done    (uSystolicPE_327_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_327_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_327_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_327_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_327_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_327_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_327_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_5_13                    ), //i
    .io_ifm_dff     (ifm_dff_x_5_13                     ), //i
    .io_wght_sign   (wght_sign_x_13_5                   ), //i
    .io_randW       (randW_x_5_13[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_13_5[14:0]              ), //i
    .io_ofm         (ofm_x_13_6[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_327_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_327_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_327_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_327_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_327_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_327_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_327_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_327_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_327_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_327_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_327_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_327_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_327_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_328 (
    .io_mac_done    (uSystolicPE_328_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_328_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_328_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_328_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_328_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_328_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_328_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_5_14                    ), //i
    .io_ifm_dff     (ifm_dff_x_5_14                     ), //i
    .io_wght_sign   (wght_sign_x_14_5                   ), //i
    .io_randW       (randW_x_5_14[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_14_5[14:0]              ), //i
    .io_ofm         (ofm_x_14_6[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_328_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_328_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_328_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_328_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_328_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_328_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_328_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_328_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_328_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_328_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_328_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_328_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_328_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_329 (
    .io_mac_done    (uSystolicPE_329_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_329_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_329_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_329_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_329_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_329_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_329_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_5_15                    ), //i
    .io_ifm_dff     (ifm_dff_x_5_15                     ), //i
    .io_wght_sign   (wght_sign_x_15_5                   ), //i
    .io_randW       (randW_x_5_15[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_15_5[14:0]              ), //i
    .io_ofm         (ofm_x_15_6[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_329_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_329_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_329_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_329_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_329_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_329_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_329_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_329_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_329_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_329_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_329_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_329_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_329_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPEBorder uSystolicPEBorder_22 (
    .io_mac_done    (uSystolicPEBorder_22_io_mac_done        ), //i
    .io_enable_i    (uSystolicPEBorder_22_io_enable_i        ), //i
    .io_clear_i     (uSystolicPEBorder_22_io_clear_i         ), //i
    .io_enable_w    (uSystolicPEBorder_22_io_enable_w        ), //i
    .io_clear_w     (uSystolicPEBorder_22_io_clear_w         ), //i
    .io_enable_o    (uSystolicPEBorder_22_io_enable_o        ), //i
    .io_clear_o     (uSystolicPEBorder_22_io_clear_o         ), //i
    .io_ifm         (io_ifm_6[15:0]                          ), //i
    .io_wght_sign   (wght_sign_x_0_6                         ), //i
    .io_wght_abs    (wght_abs_x_0_6[14:0]                    ), //i
    .io_ofm         (ofm_x_0_7[31:0]                         ), //i
    .io_mac_done_d  (uSystolicPEBorder_22_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPEBorder_22_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPEBorder_22_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPEBorder_22_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPEBorder_22_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPEBorder_22_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPEBorder_22_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPEBorder_22_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPEBorder_22_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPEBorder_22_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPEBorder_22_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPEBorder_22_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPEBorder_22_io_ofm_d[31:0]     ), //o
    .clk            (clk                                     ), //i
    .reset          (reset                                   )  //i
  );
  uSystolicPE uSystolicPE_330 (
    .io_mac_done    (uSystolicPE_330_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_330_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_330_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_330_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_330_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_330_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_330_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_6_1                     ), //i
    .io_ifm_dff     (ifm_dff_x_6_1                      ), //i
    .io_wght_sign   (wght_sign_x_1_6                    ), //i
    .io_randW       (randW_x_6_1[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_1_6[14:0]               ), //i
    .io_ofm         (ofm_x_1_7[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_330_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_330_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_330_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_330_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_330_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_330_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_330_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_330_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_330_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_330_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_330_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_330_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_330_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_331 (
    .io_mac_done    (uSystolicPE_331_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_331_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_331_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_331_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_331_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_331_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_331_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_6_2                     ), //i
    .io_ifm_dff     (ifm_dff_x_6_2                      ), //i
    .io_wght_sign   (wght_sign_x_2_6                    ), //i
    .io_randW       (randW_x_6_2[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_2_6[14:0]               ), //i
    .io_ofm         (ofm_x_2_7[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_331_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_331_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_331_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_331_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_331_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_331_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_331_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_331_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_331_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_331_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_331_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_331_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_331_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_332 (
    .io_mac_done    (uSystolicPE_332_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_332_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_332_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_332_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_332_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_332_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_332_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_6_3                     ), //i
    .io_ifm_dff     (ifm_dff_x_6_3                      ), //i
    .io_wght_sign   (wght_sign_x_3_6                    ), //i
    .io_randW       (randW_x_6_3[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_3_6[14:0]               ), //i
    .io_ofm         (ofm_x_3_7[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_332_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_332_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_332_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_332_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_332_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_332_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_332_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_332_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_332_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_332_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_332_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_332_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_332_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_333 (
    .io_mac_done    (uSystolicPE_333_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_333_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_333_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_333_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_333_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_333_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_333_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_6_4                     ), //i
    .io_ifm_dff     (ifm_dff_x_6_4                      ), //i
    .io_wght_sign   (wght_sign_x_4_6                    ), //i
    .io_randW       (randW_x_6_4[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_4_6[14:0]               ), //i
    .io_ofm         (ofm_x_4_7[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_333_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_333_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_333_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_333_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_333_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_333_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_333_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_333_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_333_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_333_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_333_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_333_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_333_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_334 (
    .io_mac_done    (uSystolicPE_334_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_334_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_334_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_334_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_334_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_334_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_334_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_6_5                     ), //i
    .io_ifm_dff     (ifm_dff_x_6_5                      ), //i
    .io_wght_sign   (wght_sign_x_5_6                    ), //i
    .io_randW       (randW_x_6_5[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_5_6[14:0]               ), //i
    .io_ofm         (ofm_x_5_7[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_334_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_334_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_334_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_334_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_334_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_334_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_334_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_334_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_334_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_334_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_334_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_334_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_334_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_335 (
    .io_mac_done    (uSystolicPE_335_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_335_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_335_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_335_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_335_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_335_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_335_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_6_6                     ), //i
    .io_ifm_dff     (ifm_dff_x_6_6                      ), //i
    .io_wght_sign   (wght_sign_x_6_6                    ), //i
    .io_randW       (randW_x_6_6[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_6_6[14:0]               ), //i
    .io_ofm         (ofm_x_6_7[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_335_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_335_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_335_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_335_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_335_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_335_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_335_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_335_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_335_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_335_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_335_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_335_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_335_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_336 (
    .io_mac_done    (uSystolicPE_336_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_336_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_336_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_336_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_336_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_336_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_336_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_6_7                     ), //i
    .io_ifm_dff     (ifm_dff_x_6_7                      ), //i
    .io_wght_sign   (wght_sign_x_7_6                    ), //i
    .io_randW       (randW_x_6_7[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_7_6[14:0]               ), //i
    .io_ofm         (ofm_x_7_7[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_336_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_336_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_336_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_336_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_336_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_336_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_336_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_336_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_336_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_336_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_336_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_336_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_336_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_337 (
    .io_mac_done    (uSystolicPE_337_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_337_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_337_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_337_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_337_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_337_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_337_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_6_8                     ), //i
    .io_ifm_dff     (ifm_dff_x_6_8                      ), //i
    .io_wght_sign   (wght_sign_x_8_6                    ), //i
    .io_randW       (randW_x_6_8[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_8_6[14:0]               ), //i
    .io_ofm         (ofm_x_8_7[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_337_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_337_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_337_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_337_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_337_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_337_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_337_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_337_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_337_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_337_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_337_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_337_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_337_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_338 (
    .io_mac_done    (uSystolicPE_338_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_338_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_338_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_338_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_338_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_338_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_338_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_6_9                     ), //i
    .io_ifm_dff     (ifm_dff_x_6_9                      ), //i
    .io_wght_sign   (wght_sign_x_9_6                    ), //i
    .io_randW       (randW_x_6_9[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_9_6[14:0]               ), //i
    .io_ofm         (ofm_x_9_7[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_338_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_338_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_338_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_338_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_338_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_338_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_338_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_338_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_338_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_338_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_338_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_338_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_338_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_339 (
    .io_mac_done    (uSystolicPE_339_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_339_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_339_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_339_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_339_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_339_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_339_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_6_10                    ), //i
    .io_ifm_dff     (ifm_dff_x_6_10                     ), //i
    .io_wght_sign   (wght_sign_x_10_6                   ), //i
    .io_randW       (randW_x_6_10[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_10_6[14:0]              ), //i
    .io_ofm         (ofm_x_10_7[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_339_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_339_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_339_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_339_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_339_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_339_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_339_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_339_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_339_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_339_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_339_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_339_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_339_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_340 (
    .io_mac_done    (uSystolicPE_340_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_340_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_340_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_340_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_340_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_340_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_340_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_6_11                    ), //i
    .io_ifm_dff     (ifm_dff_x_6_11                     ), //i
    .io_wght_sign   (wght_sign_x_11_6                   ), //i
    .io_randW       (randW_x_6_11[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_11_6[14:0]              ), //i
    .io_ofm         (ofm_x_11_7[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_340_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_340_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_340_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_340_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_340_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_340_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_340_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_340_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_340_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_340_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_340_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_340_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_340_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_341 (
    .io_mac_done    (uSystolicPE_341_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_341_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_341_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_341_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_341_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_341_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_341_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_6_12                    ), //i
    .io_ifm_dff     (ifm_dff_x_6_12                     ), //i
    .io_wght_sign   (wght_sign_x_12_6                   ), //i
    .io_randW       (randW_x_6_12[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_12_6[14:0]              ), //i
    .io_ofm         (ofm_x_12_7[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_341_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_341_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_341_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_341_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_341_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_341_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_341_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_341_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_341_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_341_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_341_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_341_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_341_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_342 (
    .io_mac_done    (uSystolicPE_342_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_342_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_342_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_342_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_342_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_342_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_342_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_6_13                    ), //i
    .io_ifm_dff     (ifm_dff_x_6_13                     ), //i
    .io_wght_sign   (wght_sign_x_13_6                   ), //i
    .io_randW       (randW_x_6_13[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_13_6[14:0]              ), //i
    .io_ofm         (ofm_x_13_7[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_342_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_342_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_342_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_342_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_342_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_342_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_342_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_342_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_342_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_342_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_342_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_342_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_342_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_343 (
    .io_mac_done    (uSystolicPE_343_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_343_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_343_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_343_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_343_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_343_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_343_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_6_14                    ), //i
    .io_ifm_dff     (ifm_dff_x_6_14                     ), //i
    .io_wght_sign   (wght_sign_x_14_6                   ), //i
    .io_randW       (randW_x_6_14[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_14_6[14:0]              ), //i
    .io_ofm         (ofm_x_14_7[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_343_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_343_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_343_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_343_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_343_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_343_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_343_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_343_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_343_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_343_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_343_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_343_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_343_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_344 (
    .io_mac_done    (uSystolicPE_344_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_344_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_344_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_344_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_344_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_344_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_344_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_6_15                    ), //i
    .io_ifm_dff     (ifm_dff_x_6_15                     ), //i
    .io_wght_sign   (wght_sign_x_15_6                   ), //i
    .io_randW       (randW_x_6_15[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_15_6[14:0]              ), //i
    .io_ofm         (ofm_x_15_7[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_344_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_344_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_344_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_344_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_344_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_344_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_344_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_344_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_344_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_344_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_344_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_344_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_344_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPEBorder uSystolicPEBorder_23 (
    .io_mac_done    (uSystolicPEBorder_23_io_mac_done        ), //i
    .io_enable_i    (uSystolicPEBorder_23_io_enable_i        ), //i
    .io_clear_i     (uSystolicPEBorder_23_io_clear_i         ), //i
    .io_enable_w    (uSystolicPEBorder_23_io_enable_w        ), //i
    .io_clear_w     (uSystolicPEBorder_23_io_clear_w         ), //i
    .io_enable_o    (uSystolicPEBorder_23_io_enable_o        ), //i
    .io_clear_o     (uSystolicPEBorder_23_io_clear_o         ), //i
    .io_ifm         (io_ifm_7[15:0]                          ), //i
    .io_wght_sign   (wght_sign_x_0_7                         ), //i
    .io_wght_abs    (wght_abs_x_0_7[14:0]                    ), //i
    .io_ofm         (ofm_x_0_8[31:0]                         ), //i
    .io_mac_done_d  (uSystolicPEBorder_23_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPEBorder_23_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPEBorder_23_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPEBorder_23_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPEBorder_23_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPEBorder_23_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPEBorder_23_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPEBorder_23_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPEBorder_23_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPEBorder_23_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPEBorder_23_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPEBorder_23_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPEBorder_23_io_ofm_d[31:0]     ), //o
    .clk            (clk                                     ), //i
    .reset          (reset                                   )  //i
  );
  uSystolicPE uSystolicPE_345 (
    .io_mac_done    (uSystolicPE_345_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_345_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_345_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_345_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_345_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_345_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_345_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_7_1                     ), //i
    .io_ifm_dff     (ifm_dff_x_7_1                      ), //i
    .io_wght_sign   (wght_sign_x_1_7                    ), //i
    .io_randW       (randW_x_7_1[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_1_7[14:0]               ), //i
    .io_ofm         (ofm_x_1_8[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_345_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_345_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_345_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_345_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_345_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_345_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_345_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_345_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_345_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_345_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_345_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_345_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_345_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_346 (
    .io_mac_done    (uSystolicPE_346_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_346_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_346_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_346_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_346_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_346_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_346_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_7_2                     ), //i
    .io_ifm_dff     (ifm_dff_x_7_2                      ), //i
    .io_wght_sign   (wght_sign_x_2_7                    ), //i
    .io_randW       (randW_x_7_2[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_2_7[14:0]               ), //i
    .io_ofm         (ofm_x_2_8[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_346_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_346_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_346_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_346_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_346_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_346_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_346_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_346_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_346_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_346_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_346_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_346_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_346_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_347 (
    .io_mac_done    (uSystolicPE_347_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_347_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_347_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_347_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_347_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_347_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_347_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_7_3                     ), //i
    .io_ifm_dff     (ifm_dff_x_7_3                      ), //i
    .io_wght_sign   (wght_sign_x_3_7                    ), //i
    .io_randW       (randW_x_7_3[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_3_7[14:0]               ), //i
    .io_ofm         (ofm_x_3_8[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_347_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_347_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_347_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_347_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_347_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_347_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_347_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_347_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_347_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_347_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_347_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_347_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_347_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_348 (
    .io_mac_done    (uSystolicPE_348_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_348_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_348_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_348_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_348_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_348_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_348_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_7_4                     ), //i
    .io_ifm_dff     (ifm_dff_x_7_4                      ), //i
    .io_wght_sign   (wght_sign_x_4_7                    ), //i
    .io_randW       (randW_x_7_4[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_4_7[14:0]               ), //i
    .io_ofm         (ofm_x_4_8[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_348_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_348_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_348_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_348_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_348_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_348_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_348_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_348_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_348_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_348_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_348_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_348_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_348_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_349 (
    .io_mac_done    (uSystolicPE_349_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_349_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_349_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_349_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_349_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_349_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_349_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_7_5                     ), //i
    .io_ifm_dff     (ifm_dff_x_7_5                      ), //i
    .io_wght_sign   (wght_sign_x_5_7                    ), //i
    .io_randW       (randW_x_7_5[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_5_7[14:0]               ), //i
    .io_ofm         (ofm_x_5_8[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_349_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_349_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_349_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_349_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_349_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_349_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_349_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_349_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_349_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_349_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_349_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_349_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_349_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_350 (
    .io_mac_done    (uSystolicPE_350_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_350_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_350_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_350_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_350_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_350_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_350_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_7_6                     ), //i
    .io_ifm_dff     (ifm_dff_x_7_6                      ), //i
    .io_wght_sign   (wght_sign_x_6_7                    ), //i
    .io_randW       (randW_x_7_6[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_6_7[14:0]               ), //i
    .io_ofm         (ofm_x_6_8[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_350_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_350_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_350_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_350_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_350_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_350_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_350_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_350_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_350_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_350_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_350_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_350_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_350_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_351 (
    .io_mac_done    (uSystolicPE_351_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_351_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_351_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_351_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_351_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_351_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_351_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_7_7                     ), //i
    .io_ifm_dff     (ifm_dff_x_7_7                      ), //i
    .io_wght_sign   (wght_sign_x_7_7                    ), //i
    .io_randW       (randW_x_7_7[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_7_7[14:0]               ), //i
    .io_ofm         (ofm_x_7_8[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_351_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_351_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_351_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_351_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_351_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_351_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_351_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_351_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_351_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_351_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_351_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_351_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_351_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_352 (
    .io_mac_done    (uSystolicPE_352_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_352_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_352_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_352_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_352_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_352_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_352_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_7_8                     ), //i
    .io_ifm_dff     (ifm_dff_x_7_8                      ), //i
    .io_wght_sign   (wght_sign_x_8_7                    ), //i
    .io_randW       (randW_x_7_8[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_8_7[14:0]               ), //i
    .io_ofm         (ofm_x_8_8[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_352_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_352_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_352_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_352_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_352_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_352_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_352_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_352_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_352_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_352_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_352_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_352_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_352_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_353 (
    .io_mac_done    (uSystolicPE_353_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_353_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_353_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_353_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_353_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_353_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_353_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_7_9                     ), //i
    .io_ifm_dff     (ifm_dff_x_7_9                      ), //i
    .io_wght_sign   (wght_sign_x_9_7                    ), //i
    .io_randW       (randW_x_7_9[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_9_7[14:0]               ), //i
    .io_ofm         (ofm_x_9_8[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_353_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_353_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_353_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_353_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_353_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_353_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_353_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_353_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_353_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_353_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_353_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_353_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_353_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_354 (
    .io_mac_done    (uSystolicPE_354_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_354_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_354_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_354_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_354_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_354_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_354_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_7_10                    ), //i
    .io_ifm_dff     (ifm_dff_x_7_10                     ), //i
    .io_wght_sign   (wght_sign_x_10_7                   ), //i
    .io_randW       (randW_x_7_10[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_10_7[14:0]              ), //i
    .io_ofm         (ofm_x_10_8[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_354_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_354_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_354_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_354_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_354_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_354_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_354_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_354_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_354_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_354_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_354_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_354_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_354_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_355 (
    .io_mac_done    (uSystolicPE_355_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_355_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_355_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_355_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_355_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_355_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_355_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_7_11                    ), //i
    .io_ifm_dff     (ifm_dff_x_7_11                     ), //i
    .io_wght_sign   (wght_sign_x_11_7                   ), //i
    .io_randW       (randW_x_7_11[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_11_7[14:0]              ), //i
    .io_ofm         (ofm_x_11_8[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_355_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_355_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_355_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_355_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_355_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_355_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_355_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_355_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_355_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_355_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_355_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_355_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_355_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_356 (
    .io_mac_done    (uSystolicPE_356_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_356_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_356_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_356_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_356_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_356_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_356_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_7_12                    ), //i
    .io_ifm_dff     (ifm_dff_x_7_12                     ), //i
    .io_wght_sign   (wght_sign_x_12_7                   ), //i
    .io_randW       (randW_x_7_12[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_12_7[14:0]              ), //i
    .io_ofm         (ofm_x_12_8[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_356_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_356_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_356_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_356_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_356_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_356_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_356_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_356_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_356_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_356_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_356_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_356_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_356_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_357 (
    .io_mac_done    (uSystolicPE_357_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_357_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_357_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_357_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_357_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_357_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_357_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_7_13                    ), //i
    .io_ifm_dff     (ifm_dff_x_7_13                     ), //i
    .io_wght_sign   (wght_sign_x_13_7                   ), //i
    .io_randW       (randW_x_7_13[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_13_7[14:0]              ), //i
    .io_ofm         (ofm_x_13_8[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_357_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_357_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_357_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_357_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_357_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_357_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_357_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_357_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_357_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_357_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_357_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_357_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_357_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_358 (
    .io_mac_done    (uSystolicPE_358_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_358_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_358_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_358_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_358_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_358_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_358_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_7_14                    ), //i
    .io_ifm_dff     (ifm_dff_x_7_14                     ), //i
    .io_wght_sign   (wght_sign_x_14_7                   ), //i
    .io_randW       (randW_x_7_14[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_14_7[14:0]              ), //i
    .io_ofm         (ofm_x_14_8[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_358_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_358_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_358_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_358_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_358_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_358_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_358_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_358_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_358_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_358_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_358_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_358_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_358_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_359 (
    .io_mac_done    (uSystolicPE_359_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_359_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_359_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_359_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_359_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_359_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_359_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_7_15                    ), //i
    .io_ifm_dff     (ifm_dff_x_7_15                     ), //i
    .io_wght_sign   (wght_sign_x_15_7                   ), //i
    .io_randW       (randW_x_7_15[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_15_7[14:0]              ), //i
    .io_ofm         (ofm_x_15_8[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_359_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_359_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_359_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_359_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_359_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_359_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_359_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_359_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_359_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_359_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_359_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_359_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_359_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPEBorder uSystolicPEBorder_24 (
    .io_mac_done    (uSystolicPEBorder_24_io_mac_done        ), //i
    .io_enable_i    (uSystolicPEBorder_24_io_enable_i        ), //i
    .io_clear_i     (uSystolicPEBorder_24_io_clear_i         ), //i
    .io_enable_w    (uSystolicPEBorder_24_io_enable_w        ), //i
    .io_clear_w     (uSystolicPEBorder_24_io_clear_w         ), //i
    .io_enable_o    (uSystolicPEBorder_24_io_enable_o        ), //i
    .io_clear_o     (uSystolicPEBorder_24_io_clear_o         ), //i
    .io_ifm         (io_ifm_8[15:0]                          ), //i
    .io_wght_sign   (wght_sign_x_0_8                         ), //i
    .io_wght_abs    (wght_abs_x_0_8[14:0]                    ), //i
    .io_ofm         (ofm_x_0_9[31:0]                         ), //i
    .io_mac_done_d  (uSystolicPEBorder_24_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPEBorder_24_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPEBorder_24_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPEBorder_24_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPEBorder_24_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPEBorder_24_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPEBorder_24_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPEBorder_24_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPEBorder_24_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPEBorder_24_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPEBorder_24_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPEBorder_24_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPEBorder_24_io_ofm_d[31:0]     ), //o
    .clk            (clk                                     ), //i
    .reset          (reset                                   )  //i
  );
  uSystolicPE uSystolicPE_360 (
    .io_mac_done    (uSystolicPE_360_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_360_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_360_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_360_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_360_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_360_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_360_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_8_1                     ), //i
    .io_ifm_dff     (ifm_dff_x_8_1                      ), //i
    .io_wght_sign   (wght_sign_x_1_8                    ), //i
    .io_randW       (randW_x_8_1[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_1_8[14:0]               ), //i
    .io_ofm         (ofm_x_1_9[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_360_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_360_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_360_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_360_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_360_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_360_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_360_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_360_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_360_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_360_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_360_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_360_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_360_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_361 (
    .io_mac_done    (uSystolicPE_361_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_361_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_361_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_361_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_361_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_361_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_361_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_8_2                     ), //i
    .io_ifm_dff     (ifm_dff_x_8_2                      ), //i
    .io_wght_sign   (wght_sign_x_2_8                    ), //i
    .io_randW       (randW_x_8_2[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_2_8[14:0]               ), //i
    .io_ofm         (ofm_x_2_9[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_361_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_361_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_361_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_361_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_361_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_361_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_361_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_361_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_361_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_361_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_361_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_361_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_361_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_362 (
    .io_mac_done    (uSystolicPE_362_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_362_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_362_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_362_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_362_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_362_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_362_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_8_3                     ), //i
    .io_ifm_dff     (ifm_dff_x_8_3                      ), //i
    .io_wght_sign   (wght_sign_x_3_8                    ), //i
    .io_randW       (randW_x_8_3[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_3_8[14:0]               ), //i
    .io_ofm         (ofm_x_3_9[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_362_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_362_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_362_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_362_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_362_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_362_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_362_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_362_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_362_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_362_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_362_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_362_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_362_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_363 (
    .io_mac_done    (uSystolicPE_363_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_363_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_363_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_363_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_363_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_363_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_363_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_8_4                     ), //i
    .io_ifm_dff     (ifm_dff_x_8_4                      ), //i
    .io_wght_sign   (wght_sign_x_4_8                    ), //i
    .io_randW       (randW_x_8_4[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_4_8[14:0]               ), //i
    .io_ofm         (ofm_x_4_9[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_363_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_363_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_363_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_363_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_363_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_363_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_363_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_363_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_363_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_363_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_363_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_363_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_363_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_364 (
    .io_mac_done    (uSystolicPE_364_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_364_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_364_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_364_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_364_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_364_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_364_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_8_5                     ), //i
    .io_ifm_dff     (ifm_dff_x_8_5                      ), //i
    .io_wght_sign   (wght_sign_x_5_8                    ), //i
    .io_randW       (randW_x_8_5[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_5_8[14:0]               ), //i
    .io_ofm         (ofm_x_5_9[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_364_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_364_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_364_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_364_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_364_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_364_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_364_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_364_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_364_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_364_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_364_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_364_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_364_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_365 (
    .io_mac_done    (uSystolicPE_365_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_365_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_365_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_365_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_365_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_365_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_365_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_8_6                     ), //i
    .io_ifm_dff     (ifm_dff_x_8_6                      ), //i
    .io_wght_sign   (wght_sign_x_6_8                    ), //i
    .io_randW       (randW_x_8_6[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_6_8[14:0]               ), //i
    .io_ofm         (ofm_x_6_9[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_365_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_365_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_365_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_365_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_365_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_365_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_365_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_365_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_365_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_365_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_365_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_365_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_365_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_366 (
    .io_mac_done    (uSystolicPE_366_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_366_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_366_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_366_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_366_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_366_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_366_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_8_7                     ), //i
    .io_ifm_dff     (ifm_dff_x_8_7                      ), //i
    .io_wght_sign   (wght_sign_x_7_8                    ), //i
    .io_randW       (randW_x_8_7[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_7_8[14:0]               ), //i
    .io_ofm         (ofm_x_7_9[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_366_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_366_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_366_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_366_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_366_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_366_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_366_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_366_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_366_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_366_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_366_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_366_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_366_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_367 (
    .io_mac_done    (uSystolicPE_367_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_367_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_367_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_367_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_367_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_367_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_367_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_8_8                     ), //i
    .io_ifm_dff     (ifm_dff_x_8_8                      ), //i
    .io_wght_sign   (wght_sign_x_8_8                    ), //i
    .io_randW       (randW_x_8_8[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_8_8[14:0]               ), //i
    .io_ofm         (ofm_x_8_9[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_367_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_367_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_367_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_367_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_367_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_367_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_367_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_367_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_367_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_367_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_367_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_367_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_367_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_368 (
    .io_mac_done    (uSystolicPE_368_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_368_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_368_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_368_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_368_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_368_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_368_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_8_9                     ), //i
    .io_ifm_dff     (ifm_dff_x_8_9                      ), //i
    .io_wght_sign   (wght_sign_x_9_8                    ), //i
    .io_randW       (randW_x_8_9[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_9_8[14:0]               ), //i
    .io_ofm         (ofm_x_9_9[31:0]                    ), //i
    .io_mac_done_d  (uSystolicPE_368_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_368_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_368_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_368_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_368_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_368_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_368_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_368_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_368_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_368_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_368_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_368_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_368_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_369 (
    .io_mac_done    (uSystolicPE_369_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_369_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_369_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_369_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_369_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_369_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_369_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_8_10                    ), //i
    .io_ifm_dff     (ifm_dff_x_8_10                     ), //i
    .io_wght_sign   (wght_sign_x_10_8                   ), //i
    .io_randW       (randW_x_8_10[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_10_8[14:0]              ), //i
    .io_ofm         (ofm_x_10_9[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_369_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_369_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_369_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_369_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_369_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_369_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_369_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_369_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_369_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_369_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_369_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_369_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_369_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_370 (
    .io_mac_done    (uSystolicPE_370_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_370_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_370_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_370_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_370_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_370_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_370_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_8_11                    ), //i
    .io_ifm_dff     (ifm_dff_x_8_11                     ), //i
    .io_wght_sign   (wght_sign_x_11_8                   ), //i
    .io_randW       (randW_x_8_11[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_11_8[14:0]              ), //i
    .io_ofm         (ofm_x_11_9[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_370_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_370_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_370_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_370_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_370_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_370_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_370_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_370_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_370_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_370_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_370_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_370_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_370_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_371 (
    .io_mac_done    (uSystolicPE_371_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_371_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_371_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_371_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_371_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_371_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_371_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_8_12                    ), //i
    .io_ifm_dff     (ifm_dff_x_8_12                     ), //i
    .io_wght_sign   (wght_sign_x_12_8                   ), //i
    .io_randW       (randW_x_8_12[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_12_8[14:0]              ), //i
    .io_ofm         (ofm_x_12_9[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_371_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_371_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_371_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_371_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_371_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_371_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_371_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_371_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_371_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_371_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_371_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_371_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_371_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_372 (
    .io_mac_done    (uSystolicPE_372_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_372_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_372_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_372_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_372_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_372_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_372_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_8_13                    ), //i
    .io_ifm_dff     (ifm_dff_x_8_13                     ), //i
    .io_wght_sign   (wght_sign_x_13_8                   ), //i
    .io_randW       (randW_x_8_13[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_13_8[14:0]              ), //i
    .io_ofm         (ofm_x_13_9[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_372_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_372_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_372_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_372_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_372_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_372_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_372_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_372_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_372_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_372_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_372_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_372_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_372_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_373 (
    .io_mac_done    (uSystolicPE_373_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_373_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_373_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_373_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_373_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_373_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_373_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_8_14                    ), //i
    .io_ifm_dff     (ifm_dff_x_8_14                     ), //i
    .io_wght_sign   (wght_sign_x_14_8                   ), //i
    .io_randW       (randW_x_8_14[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_14_8[14:0]              ), //i
    .io_ofm         (ofm_x_14_9[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_373_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_373_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_373_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_373_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_373_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_373_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_373_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_373_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_373_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_373_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_373_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_373_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_373_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_374 (
    .io_mac_done    (uSystolicPE_374_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_374_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_374_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_374_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_374_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_374_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_374_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_8_15                    ), //i
    .io_ifm_dff     (ifm_dff_x_8_15                     ), //i
    .io_wght_sign   (wght_sign_x_15_8                   ), //i
    .io_randW       (randW_x_8_15[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_15_8[14:0]              ), //i
    .io_ofm         (ofm_x_15_9[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_374_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_374_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_374_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_374_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_374_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_374_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_374_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_374_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_374_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_374_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_374_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_374_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_374_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPEBorder uSystolicPEBorder_25 (
    .io_mac_done    (uSystolicPEBorder_25_io_mac_done        ), //i
    .io_enable_i    (uSystolicPEBorder_25_io_enable_i        ), //i
    .io_clear_i     (uSystolicPEBorder_25_io_clear_i         ), //i
    .io_enable_w    (uSystolicPEBorder_25_io_enable_w        ), //i
    .io_clear_w     (uSystolicPEBorder_25_io_clear_w         ), //i
    .io_enable_o    (uSystolicPEBorder_25_io_enable_o        ), //i
    .io_clear_o     (uSystolicPEBorder_25_io_clear_o         ), //i
    .io_ifm         (io_ifm_9[15:0]                          ), //i
    .io_wght_sign   (wght_sign_x_0_9                         ), //i
    .io_wght_abs    (wght_abs_x_0_9[14:0]                    ), //i
    .io_ofm         (ofm_x_0_10[31:0]                        ), //i
    .io_mac_done_d  (uSystolicPEBorder_25_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPEBorder_25_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPEBorder_25_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPEBorder_25_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPEBorder_25_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPEBorder_25_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPEBorder_25_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPEBorder_25_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPEBorder_25_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPEBorder_25_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPEBorder_25_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPEBorder_25_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPEBorder_25_io_ofm_d[31:0]     ), //o
    .clk            (clk                                     ), //i
    .reset          (reset                                   )  //i
  );
  uSystolicPE uSystolicPE_375 (
    .io_mac_done    (uSystolicPE_375_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_375_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_375_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_375_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_375_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_375_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_375_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_9_1                     ), //i
    .io_ifm_dff     (ifm_dff_x_9_1                      ), //i
    .io_wght_sign   (wght_sign_x_1_9                    ), //i
    .io_randW       (randW_x_9_1[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_1_9[14:0]               ), //i
    .io_ofm         (ofm_x_1_10[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_375_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_375_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_375_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_375_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_375_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_375_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_375_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_375_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_375_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_375_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_375_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_375_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_375_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_376 (
    .io_mac_done    (uSystolicPE_376_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_376_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_376_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_376_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_376_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_376_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_376_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_9_2                     ), //i
    .io_ifm_dff     (ifm_dff_x_9_2                      ), //i
    .io_wght_sign   (wght_sign_x_2_9                    ), //i
    .io_randW       (randW_x_9_2[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_2_9[14:0]               ), //i
    .io_ofm         (ofm_x_2_10[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_376_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_376_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_376_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_376_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_376_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_376_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_376_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_376_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_376_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_376_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_376_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_376_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_376_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_377 (
    .io_mac_done    (uSystolicPE_377_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_377_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_377_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_377_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_377_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_377_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_377_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_9_3                     ), //i
    .io_ifm_dff     (ifm_dff_x_9_3                      ), //i
    .io_wght_sign   (wght_sign_x_3_9                    ), //i
    .io_randW       (randW_x_9_3[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_3_9[14:0]               ), //i
    .io_ofm         (ofm_x_3_10[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_377_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_377_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_377_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_377_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_377_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_377_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_377_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_377_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_377_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_377_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_377_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_377_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_377_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_378 (
    .io_mac_done    (uSystolicPE_378_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_378_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_378_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_378_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_378_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_378_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_378_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_9_4                     ), //i
    .io_ifm_dff     (ifm_dff_x_9_4                      ), //i
    .io_wght_sign   (wght_sign_x_4_9                    ), //i
    .io_randW       (randW_x_9_4[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_4_9[14:0]               ), //i
    .io_ofm         (ofm_x_4_10[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_378_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_378_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_378_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_378_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_378_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_378_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_378_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_378_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_378_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_378_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_378_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_378_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_378_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_379 (
    .io_mac_done    (uSystolicPE_379_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_379_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_379_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_379_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_379_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_379_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_379_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_9_5                     ), //i
    .io_ifm_dff     (ifm_dff_x_9_5                      ), //i
    .io_wght_sign   (wght_sign_x_5_9                    ), //i
    .io_randW       (randW_x_9_5[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_5_9[14:0]               ), //i
    .io_ofm         (ofm_x_5_10[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_379_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_379_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_379_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_379_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_379_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_379_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_379_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_379_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_379_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_379_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_379_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_379_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_379_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_380 (
    .io_mac_done    (uSystolicPE_380_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_380_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_380_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_380_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_380_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_380_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_380_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_9_6                     ), //i
    .io_ifm_dff     (ifm_dff_x_9_6                      ), //i
    .io_wght_sign   (wght_sign_x_6_9                    ), //i
    .io_randW       (randW_x_9_6[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_6_9[14:0]               ), //i
    .io_ofm         (ofm_x_6_10[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_380_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_380_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_380_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_380_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_380_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_380_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_380_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_380_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_380_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_380_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_380_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_380_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_380_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_381 (
    .io_mac_done    (uSystolicPE_381_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_381_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_381_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_381_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_381_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_381_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_381_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_9_7                     ), //i
    .io_ifm_dff     (ifm_dff_x_9_7                      ), //i
    .io_wght_sign   (wght_sign_x_7_9                    ), //i
    .io_randW       (randW_x_9_7[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_7_9[14:0]               ), //i
    .io_ofm         (ofm_x_7_10[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_381_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_381_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_381_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_381_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_381_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_381_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_381_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_381_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_381_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_381_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_381_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_381_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_381_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_382 (
    .io_mac_done    (uSystolicPE_382_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_382_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_382_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_382_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_382_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_382_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_382_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_9_8                     ), //i
    .io_ifm_dff     (ifm_dff_x_9_8                      ), //i
    .io_wght_sign   (wght_sign_x_8_9                    ), //i
    .io_randW       (randW_x_9_8[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_8_9[14:0]               ), //i
    .io_ofm         (ofm_x_8_10[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_382_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_382_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_382_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_382_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_382_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_382_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_382_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_382_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_382_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_382_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_382_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_382_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_382_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_383 (
    .io_mac_done    (uSystolicPE_383_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_383_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_383_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_383_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_383_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_383_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_383_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_9_9                     ), //i
    .io_ifm_dff     (ifm_dff_x_9_9                      ), //i
    .io_wght_sign   (wght_sign_x_9_9                    ), //i
    .io_randW       (randW_x_9_9[14:0]                  ), //i
    .io_wght_abs    (wght_abs_x_9_9[14:0]               ), //i
    .io_ofm         (ofm_x_9_10[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_383_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_383_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_383_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_383_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_383_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_383_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_383_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_383_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_383_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_383_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_383_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_383_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_383_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_384 (
    .io_mac_done    (uSystolicPE_384_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_384_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_384_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_384_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_384_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_384_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_384_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_9_10                    ), //i
    .io_ifm_dff     (ifm_dff_x_9_10                     ), //i
    .io_wght_sign   (wght_sign_x_10_9                   ), //i
    .io_randW       (randW_x_9_10[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_10_9[14:0]              ), //i
    .io_ofm         (ofm_x_10_10[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_384_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_384_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_384_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_384_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_384_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_384_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_384_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_384_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_384_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_384_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_384_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_384_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_384_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_385 (
    .io_mac_done    (uSystolicPE_385_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_385_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_385_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_385_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_385_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_385_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_385_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_9_11                    ), //i
    .io_ifm_dff     (ifm_dff_x_9_11                     ), //i
    .io_wght_sign   (wght_sign_x_11_9                   ), //i
    .io_randW       (randW_x_9_11[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_11_9[14:0]              ), //i
    .io_ofm         (ofm_x_11_10[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_385_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_385_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_385_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_385_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_385_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_385_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_385_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_385_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_385_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_385_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_385_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_385_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_385_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_386 (
    .io_mac_done    (uSystolicPE_386_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_386_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_386_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_386_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_386_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_386_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_386_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_9_12                    ), //i
    .io_ifm_dff     (ifm_dff_x_9_12                     ), //i
    .io_wght_sign   (wght_sign_x_12_9                   ), //i
    .io_randW       (randW_x_9_12[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_12_9[14:0]              ), //i
    .io_ofm         (ofm_x_12_10[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_386_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_386_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_386_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_386_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_386_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_386_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_386_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_386_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_386_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_386_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_386_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_386_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_386_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_387 (
    .io_mac_done    (uSystolicPE_387_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_387_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_387_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_387_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_387_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_387_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_387_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_9_13                    ), //i
    .io_ifm_dff     (ifm_dff_x_9_13                     ), //i
    .io_wght_sign   (wght_sign_x_13_9                   ), //i
    .io_randW       (randW_x_9_13[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_13_9[14:0]              ), //i
    .io_ofm         (ofm_x_13_10[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_387_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_387_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_387_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_387_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_387_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_387_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_387_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_387_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_387_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_387_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_387_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_387_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_387_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_388 (
    .io_mac_done    (uSystolicPE_388_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_388_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_388_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_388_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_388_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_388_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_388_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_9_14                    ), //i
    .io_ifm_dff     (ifm_dff_x_9_14                     ), //i
    .io_wght_sign   (wght_sign_x_14_9                   ), //i
    .io_randW       (randW_x_9_14[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_14_9[14:0]              ), //i
    .io_ofm         (ofm_x_14_10[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_388_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_388_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_388_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_388_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_388_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_388_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_388_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_388_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_388_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_388_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_388_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_388_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_388_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_389 (
    .io_mac_done    (uSystolicPE_389_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_389_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_389_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_389_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_389_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_389_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_389_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_9_15                    ), //i
    .io_ifm_dff     (ifm_dff_x_9_15                     ), //i
    .io_wght_sign   (wght_sign_x_15_9                   ), //i
    .io_randW       (randW_x_9_15[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_15_9[14:0]              ), //i
    .io_ofm         (ofm_x_15_10[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_389_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_389_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_389_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_389_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_389_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_389_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_389_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_389_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_389_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_389_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_389_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_389_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_389_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPEBorder uSystolicPEBorder_26 (
    .io_mac_done    (uSystolicPEBorder_26_io_mac_done        ), //i
    .io_enable_i    (uSystolicPEBorder_26_io_enable_i        ), //i
    .io_clear_i     (uSystolicPEBorder_26_io_clear_i         ), //i
    .io_enable_w    (uSystolicPEBorder_26_io_enable_w        ), //i
    .io_clear_w     (uSystolicPEBorder_26_io_clear_w         ), //i
    .io_enable_o    (uSystolicPEBorder_26_io_enable_o        ), //i
    .io_clear_o     (uSystolicPEBorder_26_io_clear_o         ), //i
    .io_ifm         (io_ifm_10[15:0]                         ), //i
    .io_wght_sign   (wght_sign_x_0_10                        ), //i
    .io_wght_abs    (wght_abs_x_0_10[14:0]                   ), //i
    .io_ofm         (ofm_x_0_11[31:0]                        ), //i
    .io_mac_done_d  (uSystolicPEBorder_26_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPEBorder_26_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPEBorder_26_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPEBorder_26_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPEBorder_26_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPEBorder_26_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPEBorder_26_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPEBorder_26_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPEBorder_26_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPEBorder_26_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPEBorder_26_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPEBorder_26_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPEBorder_26_io_ofm_d[31:0]     ), //o
    .clk            (clk                                     ), //i
    .reset          (reset                                   )  //i
  );
  uSystolicPE uSystolicPE_390 (
    .io_mac_done    (uSystolicPE_390_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_390_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_390_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_390_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_390_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_390_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_390_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_10_1                    ), //i
    .io_ifm_dff     (ifm_dff_x_10_1                     ), //i
    .io_wght_sign   (wght_sign_x_1_10                   ), //i
    .io_randW       (randW_x_10_1[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_1_10[14:0]              ), //i
    .io_ofm         (ofm_x_1_11[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_390_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_390_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_390_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_390_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_390_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_390_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_390_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_390_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_390_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_390_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_390_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_390_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_390_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_391 (
    .io_mac_done    (uSystolicPE_391_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_391_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_391_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_391_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_391_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_391_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_391_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_10_2                    ), //i
    .io_ifm_dff     (ifm_dff_x_10_2                     ), //i
    .io_wght_sign   (wght_sign_x_2_10                   ), //i
    .io_randW       (randW_x_10_2[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_2_10[14:0]              ), //i
    .io_ofm         (ofm_x_2_11[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_391_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_391_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_391_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_391_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_391_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_391_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_391_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_391_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_391_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_391_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_391_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_391_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_391_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_392 (
    .io_mac_done    (uSystolicPE_392_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_392_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_392_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_392_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_392_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_392_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_392_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_10_3                    ), //i
    .io_ifm_dff     (ifm_dff_x_10_3                     ), //i
    .io_wght_sign   (wght_sign_x_3_10                   ), //i
    .io_randW       (randW_x_10_3[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_3_10[14:0]              ), //i
    .io_ofm         (ofm_x_3_11[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_392_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_392_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_392_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_392_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_392_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_392_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_392_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_392_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_392_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_392_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_392_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_392_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_392_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_393 (
    .io_mac_done    (uSystolicPE_393_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_393_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_393_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_393_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_393_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_393_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_393_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_10_4                    ), //i
    .io_ifm_dff     (ifm_dff_x_10_4                     ), //i
    .io_wght_sign   (wght_sign_x_4_10                   ), //i
    .io_randW       (randW_x_10_4[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_4_10[14:0]              ), //i
    .io_ofm         (ofm_x_4_11[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_393_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_393_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_393_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_393_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_393_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_393_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_393_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_393_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_393_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_393_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_393_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_393_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_393_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_394 (
    .io_mac_done    (uSystolicPE_394_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_394_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_394_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_394_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_394_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_394_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_394_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_10_5                    ), //i
    .io_ifm_dff     (ifm_dff_x_10_5                     ), //i
    .io_wght_sign   (wght_sign_x_5_10                   ), //i
    .io_randW       (randW_x_10_5[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_5_10[14:0]              ), //i
    .io_ofm         (ofm_x_5_11[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_394_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_394_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_394_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_394_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_394_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_394_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_394_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_394_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_394_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_394_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_394_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_394_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_394_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_395 (
    .io_mac_done    (uSystolicPE_395_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_395_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_395_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_395_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_395_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_395_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_395_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_10_6                    ), //i
    .io_ifm_dff     (ifm_dff_x_10_6                     ), //i
    .io_wght_sign   (wght_sign_x_6_10                   ), //i
    .io_randW       (randW_x_10_6[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_6_10[14:0]              ), //i
    .io_ofm         (ofm_x_6_11[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_395_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_395_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_395_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_395_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_395_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_395_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_395_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_395_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_395_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_395_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_395_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_395_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_395_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_396 (
    .io_mac_done    (uSystolicPE_396_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_396_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_396_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_396_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_396_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_396_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_396_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_10_7                    ), //i
    .io_ifm_dff     (ifm_dff_x_10_7                     ), //i
    .io_wght_sign   (wght_sign_x_7_10                   ), //i
    .io_randW       (randW_x_10_7[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_7_10[14:0]              ), //i
    .io_ofm         (ofm_x_7_11[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_396_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_396_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_396_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_396_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_396_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_396_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_396_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_396_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_396_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_396_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_396_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_396_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_396_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_397 (
    .io_mac_done    (uSystolicPE_397_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_397_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_397_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_397_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_397_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_397_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_397_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_10_8                    ), //i
    .io_ifm_dff     (ifm_dff_x_10_8                     ), //i
    .io_wght_sign   (wght_sign_x_8_10                   ), //i
    .io_randW       (randW_x_10_8[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_8_10[14:0]              ), //i
    .io_ofm         (ofm_x_8_11[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_397_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_397_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_397_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_397_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_397_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_397_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_397_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_397_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_397_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_397_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_397_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_397_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_397_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_398 (
    .io_mac_done    (uSystolicPE_398_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_398_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_398_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_398_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_398_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_398_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_398_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_10_9                    ), //i
    .io_ifm_dff     (ifm_dff_x_10_9                     ), //i
    .io_wght_sign   (wght_sign_x_9_10                   ), //i
    .io_randW       (randW_x_10_9[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_9_10[14:0]              ), //i
    .io_ofm         (ofm_x_9_11[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_398_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_398_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_398_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_398_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_398_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_398_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_398_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_398_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_398_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_398_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_398_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_398_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_398_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_399 (
    .io_mac_done    (uSystolicPE_399_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_399_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_399_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_399_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_399_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_399_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_399_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_10_10                   ), //i
    .io_ifm_dff     (ifm_dff_x_10_10                    ), //i
    .io_wght_sign   (wght_sign_x_10_10                  ), //i
    .io_randW       (randW_x_10_10[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_10_10[14:0]             ), //i
    .io_ofm         (ofm_x_10_11[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_399_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_399_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_399_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_399_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_399_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_399_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_399_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_399_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_399_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_399_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_399_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_399_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_399_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_400 (
    .io_mac_done    (uSystolicPE_400_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_400_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_400_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_400_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_400_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_400_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_400_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_10_11                   ), //i
    .io_ifm_dff     (ifm_dff_x_10_11                    ), //i
    .io_wght_sign   (wght_sign_x_11_10                  ), //i
    .io_randW       (randW_x_10_11[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_11_10[14:0]             ), //i
    .io_ofm         (ofm_x_11_11[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_400_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_400_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_400_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_400_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_400_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_400_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_400_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_400_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_400_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_400_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_400_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_400_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_400_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_401 (
    .io_mac_done    (uSystolicPE_401_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_401_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_401_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_401_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_401_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_401_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_401_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_10_12                   ), //i
    .io_ifm_dff     (ifm_dff_x_10_12                    ), //i
    .io_wght_sign   (wght_sign_x_12_10                  ), //i
    .io_randW       (randW_x_10_12[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_12_10[14:0]             ), //i
    .io_ofm         (ofm_x_12_11[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_401_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_401_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_401_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_401_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_401_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_401_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_401_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_401_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_401_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_401_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_401_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_401_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_401_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_402 (
    .io_mac_done    (uSystolicPE_402_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_402_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_402_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_402_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_402_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_402_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_402_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_10_13                   ), //i
    .io_ifm_dff     (ifm_dff_x_10_13                    ), //i
    .io_wght_sign   (wght_sign_x_13_10                  ), //i
    .io_randW       (randW_x_10_13[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_13_10[14:0]             ), //i
    .io_ofm         (ofm_x_13_11[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_402_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_402_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_402_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_402_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_402_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_402_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_402_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_402_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_402_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_402_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_402_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_402_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_402_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_403 (
    .io_mac_done    (uSystolicPE_403_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_403_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_403_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_403_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_403_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_403_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_403_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_10_14                   ), //i
    .io_ifm_dff     (ifm_dff_x_10_14                    ), //i
    .io_wght_sign   (wght_sign_x_14_10                  ), //i
    .io_randW       (randW_x_10_14[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_14_10[14:0]             ), //i
    .io_ofm         (ofm_x_14_11[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_403_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_403_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_403_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_403_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_403_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_403_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_403_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_403_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_403_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_403_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_403_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_403_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_403_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_404 (
    .io_mac_done    (uSystolicPE_404_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_404_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_404_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_404_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_404_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_404_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_404_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_10_15                   ), //i
    .io_ifm_dff     (ifm_dff_x_10_15                    ), //i
    .io_wght_sign   (wght_sign_x_15_10                  ), //i
    .io_randW       (randW_x_10_15[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_15_10[14:0]             ), //i
    .io_ofm         (ofm_x_15_11[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_404_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_404_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_404_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_404_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_404_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_404_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_404_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_404_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_404_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_404_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_404_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_404_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_404_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPEBorder uSystolicPEBorder_27 (
    .io_mac_done    (uSystolicPEBorder_27_io_mac_done        ), //i
    .io_enable_i    (uSystolicPEBorder_27_io_enable_i        ), //i
    .io_clear_i     (uSystolicPEBorder_27_io_clear_i         ), //i
    .io_enable_w    (uSystolicPEBorder_27_io_enable_w        ), //i
    .io_clear_w     (uSystolicPEBorder_27_io_clear_w         ), //i
    .io_enable_o    (uSystolicPEBorder_27_io_enable_o        ), //i
    .io_clear_o     (uSystolicPEBorder_27_io_clear_o         ), //i
    .io_ifm         (io_ifm_11[15:0]                         ), //i
    .io_wght_sign   (wght_sign_x_0_11                        ), //i
    .io_wght_abs    (wght_abs_x_0_11[14:0]                   ), //i
    .io_ofm         (ofm_x_0_12[31:0]                        ), //i
    .io_mac_done_d  (uSystolicPEBorder_27_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPEBorder_27_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPEBorder_27_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPEBorder_27_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPEBorder_27_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPEBorder_27_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPEBorder_27_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPEBorder_27_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPEBorder_27_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPEBorder_27_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPEBorder_27_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPEBorder_27_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPEBorder_27_io_ofm_d[31:0]     ), //o
    .clk            (clk                                     ), //i
    .reset          (reset                                   )  //i
  );
  uSystolicPE uSystolicPE_405 (
    .io_mac_done    (uSystolicPE_405_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_405_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_405_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_405_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_405_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_405_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_405_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_11_1                    ), //i
    .io_ifm_dff     (ifm_dff_x_11_1                     ), //i
    .io_wght_sign   (wght_sign_x_1_11                   ), //i
    .io_randW       (randW_x_11_1[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_1_11[14:0]              ), //i
    .io_ofm         (ofm_x_1_12[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_405_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_405_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_405_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_405_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_405_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_405_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_405_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_405_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_405_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_405_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_405_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_405_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_405_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_406 (
    .io_mac_done    (uSystolicPE_406_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_406_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_406_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_406_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_406_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_406_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_406_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_11_2                    ), //i
    .io_ifm_dff     (ifm_dff_x_11_2                     ), //i
    .io_wght_sign   (wght_sign_x_2_11                   ), //i
    .io_randW       (randW_x_11_2[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_2_11[14:0]              ), //i
    .io_ofm         (ofm_x_2_12[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_406_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_406_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_406_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_406_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_406_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_406_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_406_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_406_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_406_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_406_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_406_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_406_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_406_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_407 (
    .io_mac_done    (uSystolicPE_407_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_407_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_407_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_407_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_407_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_407_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_407_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_11_3                    ), //i
    .io_ifm_dff     (ifm_dff_x_11_3                     ), //i
    .io_wght_sign   (wght_sign_x_3_11                   ), //i
    .io_randW       (randW_x_11_3[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_3_11[14:0]              ), //i
    .io_ofm         (ofm_x_3_12[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_407_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_407_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_407_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_407_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_407_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_407_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_407_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_407_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_407_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_407_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_407_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_407_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_407_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_408 (
    .io_mac_done    (uSystolicPE_408_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_408_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_408_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_408_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_408_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_408_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_408_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_11_4                    ), //i
    .io_ifm_dff     (ifm_dff_x_11_4                     ), //i
    .io_wght_sign   (wght_sign_x_4_11                   ), //i
    .io_randW       (randW_x_11_4[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_4_11[14:0]              ), //i
    .io_ofm         (ofm_x_4_12[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_408_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_408_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_408_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_408_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_408_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_408_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_408_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_408_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_408_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_408_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_408_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_408_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_408_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_409 (
    .io_mac_done    (uSystolicPE_409_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_409_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_409_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_409_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_409_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_409_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_409_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_11_5                    ), //i
    .io_ifm_dff     (ifm_dff_x_11_5                     ), //i
    .io_wght_sign   (wght_sign_x_5_11                   ), //i
    .io_randW       (randW_x_11_5[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_5_11[14:0]              ), //i
    .io_ofm         (ofm_x_5_12[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_409_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_409_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_409_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_409_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_409_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_409_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_409_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_409_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_409_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_409_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_409_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_409_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_409_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_410 (
    .io_mac_done    (uSystolicPE_410_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_410_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_410_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_410_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_410_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_410_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_410_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_11_6                    ), //i
    .io_ifm_dff     (ifm_dff_x_11_6                     ), //i
    .io_wght_sign   (wght_sign_x_6_11                   ), //i
    .io_randW       (randW_x_11_6[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_6_11[14:0]              ), //i
    .io_ofm         (ofm_x_6_12[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_410_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_410_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_410_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_410_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_410_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_410_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_410_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_410_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_410_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_410_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_410_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_410_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_410_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_411 (
    .io_mac_done    (uSystolicPE_411_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_411_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_411_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_411_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_411_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_411_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_411_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_11_7                    ), //i
    .io_ifm_dff     (ifm_dff_x_11_7                     ), //i
    .io_wght_sign   (wght_sign_x_7_11                   ), //i
    .io_randW       (randW_x_11_7[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_7_11[14:0]              ), //i
    .io_ofm         (ofm_x_7_12[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_411_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_411_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_411_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_411_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_411_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_411_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_411_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_411_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_411_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_411_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_411_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_411_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_411_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_412 (
    .io_mac_done    (uSystolicPE_412_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_412_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_412_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_412_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_412_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_412_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_412_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_11_8                    ), //i
    .io_ifm_dff     (ifm_dff_x_11_8                     ), //i
    .io_wght_sign   (wght_sign_x_8_11                   ), //i
    .io_randW       (randW_x_11_8[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_8_11[14:0]              ), //i
    .io_ofm         (ofm_x_8_12[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_412_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_412_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_412_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_412_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_412_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_412_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_412_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_412_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_412_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_412_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_412_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_412_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_412_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_413 (
    .io_mac_done    (uSystolicPE_413_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_413_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_413_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_413_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_413_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_413_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_413_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_11_9                    ), //i
    .io_ifm_dff     (ifm_dff_x_11_9                     ), //i
    .io_wght_sign   (wght_sign_x_9_11                   ), //i
    .io_randW       (randW_x_11_9[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_9_11[14:0]              ), //i
    .io_ofm         (ofm_x_9_12[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_413_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_413_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_413_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_413_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_413_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_413_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_413_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_413_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_413_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_413_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_413_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_413_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_413_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_414 (
    .io_mac_done    (uSystolicPE_414_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_414_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_414_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_414_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_414_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_414_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_414_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_11_10                   ), //i
    .io_ifm_dff     (ifm_dff_x_11_10                    ), //i
    .io_wght_sign   (wght_sign_x_10_11                  ), //i
    .io_randW       (randW_x_11_10[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_10_11[14:0]             ), //i
    .io_ofm         (ofm_x_10_12[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_414_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_414_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_414_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_414_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_414_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_414_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_414_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_414_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_414_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_414_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_414_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_414_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_414_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_415 (
    .io_mac_done    (uSystolicPE_415_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_415_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_415_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_415_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_415_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_415_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_415_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_11_11                   ), //i
    .io_ifm_dff     (ifm_dff_x_11_11                    ), //i
    .io_wght_sign   (wght_sign_x_11_11                  ), //i
    .io_randW       (randW_x_11_11[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_11_11[14:0]             ), //i
    .io_ofm         (ofm_x_11_12[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_415_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_415_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_415_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_415_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_415_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_415_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_415_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_415_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_415_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_415_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_415_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_415_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_415_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_416 (
    .io_mac_done    (uSystolicPE_416_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_416_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_416_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_416_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_416_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_416_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_416_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_11_12                   ), //i
    .io_ifm_dff     (ifm_dff_x_11_12                    ), //i
    .io_wght_sign   (wght_sign_x_12_11                  ), //i
    .io_randW       (randW_x_11_12[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_12_11[14:0]             ), //i
    .io_ofm         (ofm_x_12_12[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_416_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_416_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_416_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_416_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_416_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_416_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_416_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_416_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_416_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_416_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_416_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_416_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_416_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_417 (
    .io_mac_done    (uSystolicPE_417_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_417_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_417_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_417_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_417_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_417_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_417_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_11_13                   ), //i
    .io_ifm_dff     (ifm_dff_x_11_13                    ), //i
    .io_wght_sign   (wght_sign_x_13_11                  ), //i
    .io_randW       (randW_x_11_13[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_13_11[14:0]             ), //i
    .io_ofm         (ofm_x_13_12[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_417_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_417_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_417_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_417_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_417_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_417_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_417_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_417_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_417_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_417_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_417_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_417_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_417_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_418 (
    .io_mac_done    (uSystolicPE_418_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_418_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_418_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_418_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_418_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_418_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_418_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_11_14                   ), //i
    .io_ifm_dff     (ifm_dff_x_11_14                    ), //i
    .io_wght_sign   (wght_sign_x_14_11                  ), //i
    .io_randW       (randW_x_11_14[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_14_11[14:0]             ), //i
    .io_ofm         (ofm_x_14_12[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_418_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_418_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_418_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_418_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_418_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_418_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_418_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_418_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_418_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_418_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_418_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_418_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_418_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_419 (
    .io_mac_done    (uSystolicPE_419_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_419_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_419_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_419_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_419_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_419_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_419_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_11_15                   ), //i
    .io_ifm_dff     (ifm_dff_x_11_15                    ), //i
    .io_wght_sign   (wght_sign_x_15_11                  ), //i
    .io_randW       (randW_x_11_15[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_15_11[14:0]             ), //i
    .io_ofm         (ofm_x_15_12[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_419_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_419_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_419_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_419_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_419_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_419_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_419_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_419_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_419_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_419_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_419_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_419_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_419_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPEBorder uSystolicPEBorder_28 (
    .io_mac_done    (uSystolicPEBorder_28_io_mac_done        ), //i
    .io_enable_i    (uSystolicPEBorder_28_io_enable_i        ), //i
    .io_clear_i     (uSystolicPEBorder_28_io_clear_i         ), //i
    .io_enable_w    (uSystolicPEBorder_28_io_enable_w        ), //i
    .io_clear_w     (uSystolicPEBorder_28_io_clear_w         ), //i
    .io_enable_o    (uSystolicPEBorder_28_io_enable_o        ), //i
    .io_clear_o     (uSystolicPEBorder_28_io_clear_o         ), //i
    .io_ifm         (io_ifm_12[15:0]                         ), //i
    .io_wght_sign   (wght_sign_x_0_12                        ), //i
    .io_wght_abs    (wght_abs_x_0_12[14:0]                   ), //i
    .io_ofm         (ofm_x_0_13[31:0]                        ), //i
    .io_mac_done_d  (uSystolicPEBorder_28_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPEBorder_28_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPEBorder_28_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPEBorder_28_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPEBorder_28_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPEBorder_28_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPEBorder_28_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPEBorder_28_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPEBorder_28_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPEBorder_28_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPEBorder_28_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPEBorder_28_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPEBorder_28_io_ofm_d[31:0]     ), //o
    .clk            (clk                                     ), //i
    .reset          (reset                                   )  //i
  );
  uSystolicPE uSystolicPE_420 (
    .io_mac_done    (uSystolicPE_420_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_420_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_420_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_420_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_420_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_420_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_420_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_12_1                    ), //i
    .io_ifm_dff     (ifm_dff_x_12_1                     ), //i
    .io_wght_sign   (wght_sign_x_1_12                   ), //i
    .io_randW       (randW_x_12_1[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_1_12[14:0]              ), //i
    .io_ofm         (ofm_x_1_13[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_420_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_420_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_420_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_420_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_420_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_420_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_420_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_420_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_420_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_420_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_420_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_420_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_420_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_421 (
    .io_mac_done    (uSystolicPE_421_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_421_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_421_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_421_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_421_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_421_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_421_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_12_2                    ), //i
    .io_ifm_dff     (ifm_dff_x_12_2                     ), //i
    .io_wght_sign   (wght_sign_x_2_12                   ), //i
    .io_randW       (randW_x_12_2[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_2_12[14:0]              ), //i
    .io_ofm         (ofm_x_2_13[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_421_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_421_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_421_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_421_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_421_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_421_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_421_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_421_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_421_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_421_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_421_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_421_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_421_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_422 (
    .io_mac_done    (uSystolicPE_422_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_422_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_422_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_422_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_422_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_422_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_422_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_12_3                    ), //i
    .io_ifm_dff     (ifm_dff_x_12_3                     ), //i
    .io_wght_sign   (wght_sign_x_3_12                   ), //i
    .io_randW       (randW_x_12_3[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_3_12[14:0]              ), //i
    .io_ofm         (ofm_x_3_13[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_422_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_422_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_422_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_422_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_422_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_422_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_422_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_422_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_422_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_422_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_422_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_422_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_422_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_423 (
    .io_mac_done    (uSystolicPE_423_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_423_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_423_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_423_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_423_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_423_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_423_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_12_4                    ), //i
    .io_ifm_dff     (ifm_dff_x_12_4                     ), //i
    .io_wght_sign   (wght_sign_x_4_12                   ), //i
    .io_randW       (randW_x_12_4[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_4_12[14:0]              ), //i
    .io_ofm         (ofm_x_4_13[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_423_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_423_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_423_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_423_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_423_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_423_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_423_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_423_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_423_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_423_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_423_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_423_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_423_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_424 (
    .io_mac_done    (uSystolicPE_424_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_424_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_424_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_424_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_424_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_424_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_424_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_12_5                    ), //i
    .io_ifm_dff     (ifm_dff_x_12_5                     ), //i
    .io_wght_sign   (wght_sign_x_5_12                   ), //i
    .io_randW       (randW_x_12_5[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_5_12[14:0]              ), //i
    .io_ofm         (ofm_x_5_13[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_424_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_424_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_424_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_424_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_424_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_424_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_424_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_424_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_424_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_424_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_424_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_424_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_424_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_425 (
    .io_mac_done    (uSystolicPE_425_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_425_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_425_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_425_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_425_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_425_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_425_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_12_6                    ), //i
    .io_ifm_dff     (ifm_dff_x_12_6                     ), //i
    .io_wght_sign   (wght_sign_x_6_12                   ), //i
    .io_randW       (randW_x_12_6[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_6_12[14:0]              ), //i
    .io_ofm         (ofm_x_6_13[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_425_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_425_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_425_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_425_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_425_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_425_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_425_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_425_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_425_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_425_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_425_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_425_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_425_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_426 (
    .io_mac_done    (uSystolicPE_426_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_426_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_426_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_426_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_426_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_426_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_426_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_12_7                    ), //i
    .io_ifm_dff     (ifm_dff_x_12_7                     ), //i
    .io_wght_sign   (wght_sign_x_7_12                   ), //i
    .io_randW       (randW_x_12_7[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_7_12[14:0]              ), //i
    .io_ofm         (ofm_x_7_13[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_426_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_426_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_426_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_426_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_426_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_426_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_426_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_426_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_426_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_426_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_426_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_426_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_426_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_427 (
    .io_mac_done    (uSystolicPE_427_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_427_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_427_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_427_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_427_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_427_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_427_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_12_8                    ), //i
    .io_ifm_dff     (ifm_dff_x_12_8                     ), //i
    .io_wght_sign   (wght_sign_x_8_12                   ), //i
    .io_randW       (randW_x_12_8[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_8_12[14:0]              ), //i
    .io_ofm         (ofm_x_8_13[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_427_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_427_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_427_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_427_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_427_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_427_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_427_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_427_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_427_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_427_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_427_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_427_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_427_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_428 (
    .io_mac_done    (uSystolicPE_428_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_428_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_428_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_428_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_428_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_428_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_428_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_12_9                    ), //i
    .io_ifm_dff     (ifm_dff_x_12_9                     ), //i
    .io_wght_sign   (wght_sign_x_9_12                   ), //i
    .io_randW       (randW_x_12_9[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_9_12[14:0]              ), //i
    .io_ofm         (ofm_x_9_13[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_428_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_428_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_428_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_428_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_428_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_428_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_428_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_428_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_428_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_428_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_428_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_428_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_428_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_429 (
    .io_mac_done    (uSystolicPE_429_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_429_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_429_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_429_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_429_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_429_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_429_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_12_10                   ), //i
    .io_ifm_dff     (ifm_dff_x_12_10                    ), //i
    .io_wght_sign   (wght_sign_x_10_12                  ), //i
    .io_randW       (randW_x_12_10[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_10_12[14:0]             ), //i
    .io_ofm         (ofm_x_10_13[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_429_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_429_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_429_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_429_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_429_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_429_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_429_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_429_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_429_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_429_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_429_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_429_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_429_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_430 (
    .io_mac_done    (uSystolicPE_430_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_430_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_430_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_430_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_430_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_430_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_430_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_12_11                   ), //i
    .io_ifm_dff     (ifm_dff_x_12_11                    ), //i
    .io_wght_sign   (wght_sign_x_11_12                  ), //i
    .io_randW       (randW_x_12_11[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_11_12[14:0]             ), //i
    .io_ofm         (ofm_x_11_13[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_430_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_430_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_430_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_430_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_430_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_430_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_430_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_430_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_430_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_430_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_430_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_430_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_430_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_431 (
    .io_mac_done    (uSystolicPE_431_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_431_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_431_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_431_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_431_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_431_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_431_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_12_12                   ), //i
    .io_ifm_dff     (ifm_dff_x_12_12                    ), //i
    .io_wght_sign   (wght_sign_x_12_12                  ), //i
    .io_randW       (randW_x_12_12[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_12_12[14:0]             ), //i
    .io_ofm         (ofm_x_12_13[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_431_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_431_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_431_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_431_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_431_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_431_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_431_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_431_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_431_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_431_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_431_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_431_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_431_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_432 (
    .io_mac_done    (uSystolicPE_432_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_432_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_432_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_432_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_432_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_432_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_432_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_12_13                   ), //i
    .io_ifm_dff     (ifm_dff_x_12_13                    ), //i
    .io_wght_sign   (wght_sign_x_13_12                  ), //i
    .io_randW       (randW_x_12_13[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_13_12[14:0]             ), //i
    .io_ofm         (ofm_x_13_13[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_432_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_432_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_432_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_432_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_432_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_432_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_432_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_432_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_432_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_432_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_432_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_432_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_432_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_433 (
    .io_mac_done    (uSystolicPE_433_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_433_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_433_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_433_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_433_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_433_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_433_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_12_14                   ), //i
    .io_ifm_dff     (ifm_dff_x_12_14                    ), //i
    .io_wght_sign   (wght_sign_x_14_12                  ), //i
    .io_randW       (randW_x_12_14[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_14_12[14:0]             ), //i
    .io_ofm         (ofm_x_14_13[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_433_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_433_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_433_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_433_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_433_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_433_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_433_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_433_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_433_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_433_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_433_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_433_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_433_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_434 (
    .io_mac_done    (uSystolicPE_434_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_434_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_434_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_434_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_434_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_434_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_434_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_12_15                   ), //i
    .io_ifm_dff     (ifm_dff_x_12_15                    ), //i
    .io_wght_sign   (wght_sign_x_15_12                  ), //i
    .io_randW       (randW_x_12_15[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_15_12[14:0]             ), //i
    .io_ofm         (ofm_x_15_13[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_434_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_434_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_434_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_434_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_434_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_434_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_434_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_434_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_434_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_434_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_434_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_434_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_434_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPEBorder uSystolicPEBorder_29 (
    .io_mac_done    (uSystolicPEBorder_29_io_mac_done        ), //i
    .io_enable_i    (uSystolicPEBorder_29_io_enable_i        ), //i
    .io_clear_i     (uSystolicPEBorder_29_io_clear_i         ), //i
    .io_enable_w    (uSystolicPEBorder_29_io_enable_w        ), //i
    .io_clear_w     (uSystolicPEBorder_29_io_clear_w         ), //i
    .io_enable_o    (uSystolicPEBorder_29_io_enable_o        ), //i
    .io_clear_o     (uSystolicPEBorder_29_io_clear_o         ), //i
    .io_ifm         (io_ifm_13[15:0]                         ), //i
    .io_wght_sign   (wght_sign_x_0_13                        ), //i
    .io_wght_abs    (wght_abs_x_0_13[14:0]                   ), //i
    .io_ofm         (ofm_x_0_14[31:0]                        ), //i
    .io_mac_done_d  (uSystolicPEBorder_29_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPEBorder_29_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPEBorder_29_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPEBorder_29_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPEBorder_29_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPEBorder_29_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPEBorder_29_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPEBorder_29_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPEBorder_29_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPEBorder_29_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPEBorder_29_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPEBorder_29_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPEBorder_29_io_ofm_d[31:0]     ), //o
    .clk            (clk                                     ), //i
    .reset          (reset                                   )  //i
  );
  uSystolicPE uSystolicPE_435 (
    .io_mac_done    (uSystolicPE_435_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_435_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_435_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_435_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_435_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_435_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_435_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_13_1                    ), //i
    .io_ifm_dff     (ifm_dff_x_13_1                     ), //i
    .io_wght_sign   (wght_sign_x_1_13                   ), //i
    .io_randW       (randW_x_13_1[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_1_13[14:0]              ), //i
    .io_ofm         (ofm_x_1_14[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_435_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_435_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_435_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_435_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_435_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_435_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_435_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_435_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_435_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_435_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_435_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_435_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_435_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_436 (
    .io_mac_done    (uSystolicPE_436_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_436_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_436_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_436_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_436_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_436_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_436_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_13_2                    ), //i
    .io_ifm_dff     (ifm_dff_x_13_2                     ), //i
    .io_wght_sign   (wght_sign_x_2_13                   ), //i
    .io_randW       (randW_x_13_2[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_2_13[14:0]              ), //i
    .io_ofm         (ofm_x_2_14[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_436_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_436_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_436_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_436_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_436_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_436_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_436_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_436_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_436_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_436_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_436_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_436_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_436_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_437 (
    .io_mac_done    (uSystolicPE_437_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_437_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_437_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_437_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_437_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_437_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_437_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_13_3                    ), //i
    .io_ifm_dff     (ifm_dff_x_13_3                     ), //i
    .io_wght_sign   (wght_sign_x_3_13                   ), //i
    .io_randW       (randW_x_13_3[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_3_13[14:0]              ), //i
    .io_ofm         (ofm_x_3_14[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_437_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_437_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_437_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_437_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_437_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_437_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_437_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_437_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_437_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_437_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_437_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_437_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_437_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_438 (
    .io_mac_done    (uSystolicPE_438_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_438_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_438_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_438_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_438_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_438_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_438_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_13_4                    ), //i
    .io_ifm_dff     (ifm_dff_x_13_4                     ), //i
    .io_wght_sign   (wght_sign_x_4_13                   ), //i
    .io_randW       (randW_x_13_4[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_4_13[14:0]              ), //i
    .io_ofm         (ofm_x_4_14[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_438_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_438_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_438_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_438_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_438_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_438_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_438_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_438_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_438_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_438_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_438_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_438_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_438_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_439 (
    .io_mac_done    (uSystolicPE_439_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_439_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_439_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_439_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_439_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_439_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_439_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_13_5                    ), //i
    .io_ifm_dff     (ifm_dff_x_13_5                     ), //i
    .io_wght_sign   (wght_sign_x_5_13                   ), //i
    .io_randW       (randW_x_13_5[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_5_13[14:0]              ), //i
    .io_ofm         (ofm_x_5_14[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_439_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_439_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_439_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_439_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_439_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_439_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_439_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_439_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_439_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_439_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_439_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_439_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_439_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_440 (
    .io_mac_done    (uSystolicPE_440_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_440_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_440_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_440_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_440_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_440_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_440_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_13_6                    ), //i
    .io_ifm_dff     (ifm_dff_x_13_6                     ), //i
    .io_wght_sign   (wght_sign_x_6_13                   ), //i
    .io_randW       (randW_x_13_6[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_6_13[14:0]              ), //i
    .io_ofm         (ofm_x_6_14[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_440_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_440_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_440_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_440_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_440_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_440_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_440_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_440_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_440_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_440_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_440_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_440_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_440_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_441 (
    .io_mac_done    (uSystolicPE_441_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_441_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_441_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_441_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_441_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_441_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_441_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_13_7                    ), //i
    .io_ifm_dff     (ifm_dff_x_13_7                     ), //i
    .io_wght_sign   (wght_sign_x_7_13                   ), //i
    .io_randW       (randW_x_13_7[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_7_13[14:0]              ), //i
    .io_ofm         (ofm_x_7_14[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_441_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_441_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_441_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_441_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_441_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_441_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_441_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_441_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_441_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_441_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_441_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_441_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_441_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_442 (
    .io_mac_done    (uSystolicPE_442_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_442_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_442_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_442_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_442_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_442_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_442_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_13_8                    ), //i
    .io_ifm_dff     (ifm_dff_x_13_8                     ), //i
    .io_wght_sign   (wght_sign_x_8_13                   ), //i
    .io_randW       (randW_x_13_8[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_8_13[14:0]              ), //i
    .io_ofm         (ofm_x_8_14[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_442_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_442_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_442_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_442_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_442_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_442_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_442_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_442_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_442_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_442_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_442_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_442_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_442_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_443 (
    .io_mac_done    (uSystolicPE_443_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_443_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_443_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_443_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_443_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_443_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_443_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_13_9                    ), //i
    .io_ifm_dff     (ifm_dff_x_13_9                     ), //i
    .io_wght_sign   (wght_sign_x_9_13                   ), //i
    .io_randW       (randW_x_13_9[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_9_13[14:0]              ), //i
    .io_ofm         (ofm_x_9_14[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_443_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_443_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_443_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_443_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_443_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_443_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_443_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_443_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_443_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_443_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_443_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_443_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_443_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_444 (
    .io_mac_done    (uSystolicPE_444_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_444_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_444_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_444_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_444_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_444_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_444_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_13_10                   ), //i
    .io_ifm_dff     (ifm_dff_x_13_10                    ), //i
    .io_wght_sign   (wght_sign_x_10_13                  ), //i
    .io_randW       (randW_x_13_10[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_10_13[14:0]             ), //i
    .io_ofm         (ofm_x_10_14[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_444_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_444_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_444_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_444_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_444_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_444_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_444_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_444_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_444_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_444_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_444_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_444_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_444_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_445 (
    .io_mac_done    (uSystolicPE_445_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_445_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_445_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_445_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_445_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_445_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_445_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_13_11                   ), //i
    .io_ifm_dff     (ifm_dff_x_13_11                    ), //i
    .io_wght_sign   (wght_sign_x_11_13                  ), //i
    .io_randW       (randW_x_13_11[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_11_13[14:0]             ), //i
    .io_ofm         (ofm_x_11_14[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_445_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_445_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_445_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_445_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_445_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_445_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_445_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_445_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_445_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_445_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_445_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_445_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_445_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_446 (
    .io_mac_done    (uSystolicPE_446_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_446_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_446_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_446_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_446_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_446_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_446_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_13_12                   ), //i
    .io_ifm_dff     (ifm_dff_x_13_12                    ), //i
    .io_wght_sign   (wght_sign_x_12_13                  ), //i
    .io_randW       (randW_x_13_12[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_12_13[14:0]             ), //i
    .io_ofm         (ofm_x_12_14[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_446_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_446_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_446_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_446_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_446_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_446_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_446_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_446_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_446_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_446_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_446_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_446_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_446_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_447 (
    .io_mac_done    (uSystolicPE_447_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_447_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_447_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_447_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_447_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_447_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_447_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_13_13                   ), //i
    .io_ifm_dff     (ifm_dff_x_13_13                    ), //i
    .io_wght_sign   (wght_sign_x_13_13                  ), //i
    .io_randW       (randW_x_13_13[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_13_13[14:0]             ), //i
    .io_ofm         (ofm_x_13_14[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_447_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_447_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_447_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_447_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_447_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_447_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_447_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_447_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_447_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_447_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_447_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_447_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_447_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_448 (
    .io_mac_done    (uSystolicPE_448_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_448_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_448_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_448_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_448_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_448_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_448_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_13_14                   ), //i
    .io_ifm_dff     (ifm_dff_x_13_14                    ), //i
    .io_wght_sign   (wght_sign_x_14_13                  ), //i
    .io_randW       (randW_x_13_14[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_14_13[14:0]             ), //i
    .io_ofm         (ofm_x_14_14[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_448_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_448_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_448_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_448_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_448_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_448_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_448_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_448_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_448_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_448_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_448_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_448_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_448_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_449 (
    .io_mac_done    (uSystolicPE_449_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_449_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_449_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_449_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_449_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_449_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_449_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_13_15                   ), //i
    .io_ifm_dff     (ifm_dff_x_13_15                    ), //i
    .io_wght_sign   (wght_sign_x_15_13                  ), //i
    .io_randW       (randW_x_13_15[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_15_13[14:0]             ), //i
    .io_ofm         (ofm_x_15_14[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_449_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_449_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_449_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_449_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_449_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_449_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_449_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_449_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_449_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_449_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_449_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_449_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_449_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPEBorder uSystolicPEBorder_30 (
    .io_mac_done    (uSystolicPEBorder_30_io_mac_done        ), //i
    .io_enable_i    (uSystolicPEBorder_30_io_enable_i        ), //i
    .io_clear_i     (uSystolicPEBorder_30_io_clear_i         ), //i
    .io_enable_w    (uSystolicPEBorder_30_io_enable_w        ), //i
    .io_clear_w     (uSystolicPEBorder_30_io_clear_w         ), //i
    .io_enable_o    (uSystolicPEBorder_30_io_enable_o        ), //i
    .io_clear_o     (uSystolicPEBorder_30_io_clear_o         ), //i
    .io_ifm         (io_ifm_14[15:0]                         ), //i
    .io_wght_sign   (wght_sign_x_0_14                        ), //i
    .io_wght_abs    (wght_abs_x_0_14[14:0]                   ), //i
    .io_ofm         (ofm_x_0_15[31:0]                        ), //i
    .io_mac_done_d  (uSystolicPEBorder_30_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPEBorder_30_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPEBorder_30_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPEBorder_30_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPEBorder_30_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPEBorder_30_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPEBorder_30_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPEBorder_30_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPEBorder_30_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPEBorder_30_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPEBorder_30_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPEBorder_30_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPEBorder_30_io_ofm_d[31:0]     ), //o
    .clk            (clk                                     ), //i
    .reset          (reset                                   )  //i
  );
  uSystolicPE uSystolicPE_450 (
    .io_mac_done    (uSystolicPE_450_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_450_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_450_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_450_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_450_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_450_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_450_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_14_1                    ), //i
    .io_ifm_dff     (ifm_dff_x_14_1                     ), //i
    .io_wght_sign   (wght_sign_x_1_14                   ), //i
    .io_randW       (randW_x_14_1[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_1_14[14:0]              ), //i
    .io_ofm         (ofm_x_1_15[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_450_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_450_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_450_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_450_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_450_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_450_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_450_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_450_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_450_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_450_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_450_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_450_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_450_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_451 (
    .io_mac_done    (uSystolicPE_451_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_451_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_451_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_451_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_451_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_451_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_451_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_14_2                    ), //i
    .io_ifm_dff     (ifm_dff_x_14_2                     ), //i
    .io_wght_sign   (wght_sign_x_2_14                   ), //i
    .io_randW       (randW_x_14_2[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_2_14[14:0]              ), //i
    .io_ofm         (ofm_x_2_15[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_451_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_451_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_451_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_451_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_451_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_451_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_451_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_451_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_451_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_451_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_451_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_451_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_451_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_452 (
    .io_mac_done    (uSystolicPE_452_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_452_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_452_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_452_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_452_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_452_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_452_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_14_3                    ), //i
    .io_ifm_dff     (ifm_dff_x_14_3                     ), //i
    .io_wght_sign   (wght_sign_x_3_14                   ), //i
    .io_randW       (randW_x_14_3[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_3_14[14:0]              ), //i
    .io_ofm         (ofm_x_3_15[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_452_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_452_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_452_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_452_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_452_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_452_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_452_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_452_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_452_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_452_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_452_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_452_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_452_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_453 (
    .io_mac_done    (uSystolicPE_453_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_453_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_453_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_453_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_453_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_453_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_453_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_14_4                    ), //i
    .io_ifm_dff     (ifm_dff_x_14_4                     ), //i
    .io_wght_sign   (wght_sign_x_4_14                   ), //i
    .io_randW       (randW_x_14_4[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_4_14[14:0]              ), //i
    .io_ofm         (ofm_x_4_15[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_453_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_453_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_453_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_453_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_453_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_453_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_453_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_453_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_453_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_453_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_453_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_453_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_453_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_454 (
    .io_mac_done    (uSystolicPE_454_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_454_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_454_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_454_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_454_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_454_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_454_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_14_5                    ), //i
    .io_ifm_dff     (ifm_dff_x_14_5                     ), //i
    .io_wght_sign   (wght_sign_x_5_14                   ), //i
    .io_randW       (randW_x_14_5[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_5_14[14:0]              ), //i
    .io_ofm         (ofm_x_5_15[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_454_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_454_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_454_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_454_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_454_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_454_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_454_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_454_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_454_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_454_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_454_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_454_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_454_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_455 (
    .io_mac_done    (uSystolicPE_455_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_455_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_455_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_455_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_455_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_455_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_455_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_14_6                    ), //i
    .io_ifm_dff     (ifm_dff_x_14_6                     ), //i
    .io_wght_sign   (wght_sign_x_6_14                   ), //i
    .io_randW       (randW_x_14_6[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_6_14[14:0]              ), //i
    .io_ofm         (ofm_x_6_15[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_455_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_455_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_455_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_455_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_455_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_455_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_455_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_455_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_455_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_455_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_455_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_455_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_455_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_456 (
    .io_mac_done    (uSystolicPE_456_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_456_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_456_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_456_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_456_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_456_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_456_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_14_7                    ), //i
    .io_ifm_dff     (ifm_dff_x_14_7                     ), //i
    .io_wght_sign   (wght_sign_x_7_14                   ), //i
    .io_randW       (randW_x_14_7[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_7_14[14:0]              ), //i
    .io_ofm         (ofm_x_7_15[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_456_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_456_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_456_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_456_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_456_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_456_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_456_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_456_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_456_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_456_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_456_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_456_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_456_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_457 (
    .io_mac_done    (uSystolicPE_457_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_457_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_457_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_457_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_457_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_457_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_457_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_14_8                    ), //i
    .io_ifm_dff     (ifm_dff_x_14_8                     ), //i
    .io_wght_sign   (wght_sign_x_8_14                   ), //i
    .io_randW       (randW_x_14_8[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_8_14[14:0]              ), //i
    .io_ofm         (ofm_x_8_15[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_457_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_457_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_457_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_457_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_457_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_457_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_457_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_457_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_457_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_457_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_457_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_457_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_457_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_458 (
    .io_mac_done    (uSystolicPE_458_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_458_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_458_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_458_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_458_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_458_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_458_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_14_9                    ), //i
    .io_ifm_dff     (ifm_dff_x_14_9                     ), //i
    .io_wght_sign   (wght_sign_x_9_14                   ), //i
    .io_randW       (randW_x_14_9[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_9_14[14:0]              ), //i
    .io_ofm         (ofm_x_9_15[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_458_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_458_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_458_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_458_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_458_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_458_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_458_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_458_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_458_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_458_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_458_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_458_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_458_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_459 (
    .io_mac_done    (uSystolicPE_459_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_459_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_459_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_459_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_459_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_459_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_459_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_14_10                   ), //i
    .io_ifm_dff     (ifm_dff_x_14_10                    ), //i
    .io_wght_sign   (wght_sign_x_10_14                  ), //i
    .io_randW       (randW_x_14_10[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_10_14[14:0]             ), //i
    .io_ofm         (ofm_x_10_15[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_459_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_459_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_459_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_459_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_459_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_459_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_459_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_459_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_459_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_459_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_459_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_459_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_459_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_460 (
    .io_mac_done    (uSystolicPE_460_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_460_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_460_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_460_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_460_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_460_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_460_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_14_11                   ), //i
    .io_ifm_dff     (ifm_dff_x_14_11                    ), //i
    .io_wght_sign   (wght_sign_x_11_14                  ), //i
    .io_randW       (randW_x_14_11[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_11_14[14:0]             ), //i
    .io_ofm         (ofm_x_11_15[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_460_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_460_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_460_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_460_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_460_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_460_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_460_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_460_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_460_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_460_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_460_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_460_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_460_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_461 (
    .io_mac_done    (uSystolicPE_461_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_461_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_461_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_461_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_461_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_461_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_461_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_14_12                   ), //i
    .io_ifm_dff     (ifm_dff_x_14_12                    ), //i
    .io_wght_sign   (wght_sign_x_12_14                  ), //i
    .io_randW       (randW_x_14_12[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_12_14[14:0]             ), //i
    .io_ofm         (ofm_x_12_15[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_461_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_461_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_461_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_461_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_461_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_461_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_461_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_461_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_461_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_461_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_461_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_461_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_461_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_462 (
    .io_mac_done    (uSystolicPE_462_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_462_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_462_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_462_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_462_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_462_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_462_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_14_13                   ), //i
    .io_ifm_dff     (ifm_dff_x_14_13                    ), //i
    .io_wght_sign   (wght_sign_x_13_14                  ), //i
    .io_randW       (randW_x_14_13[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_13_14[14:0]             ), //i
    .io_ofm         (ofm_x_13_15[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_462_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_462_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_462_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_462_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_462_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_462_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_462_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_462_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_462_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_462_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_462_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_462_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_462_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_463 (
    .io_mac_done    (uSystolicPE_463_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_463_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_463_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_463_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_463_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_463_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_463_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_14_14                   ), //i
    .io_ifm_dff     (ifm_dff_x_14_14                    ), //i
    .io_wght_sign   (wght_sign_x_14_14                  ), //i
    .io_randW       (randW_x_14_14[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_14_14[14:0]             ), //i
    .io_ofm         (ofm_x_14_15[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_463_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_463_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_463_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_463_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_463_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_463_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_463_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_463_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_463_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_463_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_463_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_463_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_463_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_464 (
    .io_mac_done    (uSystolicPE_464_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_464_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_464_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_464_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_464_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_464_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_464_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_14_15                   ), //i
    .io_ifm_dff     (ifm_dff_x_14_15                    ), //i
    .io_wght_sign   (wght_sign_x_15_14                  ), //i
    .io_randW       (randW_x_14_15[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_15_14[14:0]             ), //i
    .io_ofm         (ofm_x_15_15[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_464_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_464_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_464_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_464_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_464_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_464_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_464_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_464_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_464_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_464_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_464_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_464_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_464_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPEBorder uSystolicPEBorder_31 (
    .io_mac_done    (uSystolicPEBorder_31_io_mac_done        ), //i
    .io_enable_i    (uSystolicPEBorder_31_io_enable_i        ), //i
    .io_clear_i     (uSystolicPEBorder_31_io_clear_i         ), //i
    .io_enable_w    (uSystolicPEBorder_31_io_enable_w        ), //i
    .io_clear_w     (uSystolicPEBorder_31_io_clear_w         ), //i
    .io_enable_o    (uSystolicPEBorder_31_io_enable_o        ), //i
    .io_clear_o     (uSystolicPEBorder_31_io_clear_o         ), //i
    .io_ifm         (io_ifm_15[15:0]                         ), //i
    .io_wght_sign   (wght_sign_x_0_15                        ), //i
    .io_wght_abs    (wght_abs_x_0_15[14:0]                   ), //i
    .io_ofm         (ofm_x_0_16[31:0]                        ), //i
    .io_mac_done_d  (uSystolicPEBorder_31_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPEBorder_31_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPEBorder_31_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPEBorder_31_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPEBorder_31_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPEBorder_31_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPEBorder_31_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPEBorder_31_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPEBorder_31_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPEBorder_31_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPEBorder_31_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPEBorder_31_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPEBorder_31_io_ofm_d[31:0]     ), //o
    .clk            (clk                                     ), //i
    .reset          (reset                                   )  //i
  );
  uSystolicPE uSystolicPE_465 (
    .io_mac_done    (uSystolicPE_465_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_465_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_465_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_465_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_465_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_465_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_465_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_15_1                    ), //i
    .io_ifm_dff     (ifm_dff_x_15_1                     ), //i
    .io_wght_sign   (wght_sign_x_1_15                   ), //i
    .io_randW       (randW_x_15_1[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_1_15[14:0]              ), //i
    .io_ofm         (ofm_x_1_16[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_465_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_465_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_465_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_465_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_465_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_465_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_465_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_465_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_465_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_465_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_465_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_465_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_465_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_466 (
    .io_mac_done    (uSystolicPE_466_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_466_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_466_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_466_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_466_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_466_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_466_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_15_2                    ), //i
    .io_ifm_dff     (ifm_dff_x_15_2                     ), //i
    .io_wght_sign   (wght_sign_x_2_15                   ), //i
    .io_randW       (randW_x_15_2[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_2_15[14:0]              ), //i
    .io_ofm         (ofm_x_2_16[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_466_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_466_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_466_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_466_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_466_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_466_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_466_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_466_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_466_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_466_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_466_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_466_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_466_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_467 (
    .io_mac_done    (uSystolicPE_467_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_467_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_467_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_467_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_467_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_467_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_467_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_15_3                    ), //i
    .io_ifm_dff     (ifm_dff_x_15_3                     ), //i
    .io_wght_sign   (wght_sign_x_3_15                   ), //i
    .io_randW       (randW_x_15_3[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_3_15[14:0]              ), //i
    .io_ofm         (ofm_x_3_16[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_467_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_467_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_467_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_467_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_467_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_467_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_467_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_467_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_467_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_467_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_467_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_467_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_467_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_468 (
    .io_mac_done    (uSystolicPE_468_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_468_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_468_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_468_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_468_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_468_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_468_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_15_4                    ), //i
    .io_ifm_dff     (ifm_dff_x_15_4                     ), //i
    .io_wght_sign   (wght_sign_x_4_15                   ), //i
    .io_randW       (randW_x_15_4[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_4_15[14:0]              ), //i
    .io_ofm         (ofm_x_4_16[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_468_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_468_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_468_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_468_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_468_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_468_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_468_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_468_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_468_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_468_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_468_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_468_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_468_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_469 (
    .io_mac_done    (uSystolicPE_469_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_469_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_469_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_469_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_469_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_469_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_469_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_15_5                    ), //i
    .io_ifm_dff     (ifm_dff_x_15_5                     ), //i
    .io_wght_sign   (wght_sign_x_5_15                   ), //i
    .io_randW       (randW_x_15_5[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_5_15[14:0]              ), //i
    .io_ofm         (ofm_x_5_16[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_469_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_469_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_469_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_469_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_469_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_469_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_469_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_469_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_469_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_469_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_469_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_469_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_469_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_470 (
    .io_mac_done    (uSystolicPE_470_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_470_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_470_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_470_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_470_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_470_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_470_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_15_6                    ), //i
    .io_ifm_dff     (ifm_dff_x_15_6                     ), //i
    .io_wght_sign   (wght_sign_x_6_15                   ), //i
    .io_randW       (randW_x_15_6[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_6_15[14:0]              ), //i
    .io_ofm         (ofm_x_6_16[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_470_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_470_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_470_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_470_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_470_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_470_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_470_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_470_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_470_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_470_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_470_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_470_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_470_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_471 (
    .io_mac_done    (uSystolicPE_471_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_471_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_471_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_471_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_471_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_471_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_471_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_15_7                    ), //i
    .io_ifm_dff     (ifm_dff_x_15_7                     ), //i
    .io_wght_sign   (wght_sign_x_7_15                   ), //i
    .io_randW       (randW_x_15_7[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_7_15[14:0]              ), //i
    .io_ofm         (ofm_x_7_16[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_471_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_471_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_471_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_471_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_471_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_471_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_471_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_471_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_471_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_471_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_471_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_471_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_471_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_472 (
    .io_mac_done    (uSystolicPE_472_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_472_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_472_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_472_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_472_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_472_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_472_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_15_8                    ), //i
    .io_ifm_dff     (ifm_dff_x_15_8                     ), //i
    .io_wght_sign   (wght_sign_x_8_15                   ), //i
    .io_randW       (randW_x_15_8[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_8_15[14:0]              ), //i
    .io_ofm         (ofm_x_8_16[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_472_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_472_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_472_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_472_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_472_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_472_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_472_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_472_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_472_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_472_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_472_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_472_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_472_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_473 (
    .io_mac_done    (uSystolicPE_473_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_473_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_473_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_473_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_473_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_473_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_473_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_15_9                    ), //i
    .io_ifm_dff     (ifm_dff_x_15_9                     ), //i
    .io_wght_sign   (wght_sign_x_9_15                   ), //i
    .io_randW       (randW_x_15_9[14:0]                 ), //i
    .io_wght_abs    (wght_abs_x_9_15[14:0]              ), //i
    .io_ofm         (ofm_x_9_16[31:0]                   ), //i
    .io_mac_done_d  (uSystolicPE_473_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_473_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_473_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_473_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_473_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_473_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_473_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_473_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_473_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_473_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_473_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_473_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_473_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_474 (
    .io_mac_done    (uSystolicPE_474_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_474_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_474_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_474_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_474_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_474_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_474_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_15_10                   ), //i
    .io_ifm_dff     (ifm_dff_x_15_10                    ), //i
    .io_wght_sign   (wght_sign_x_10_15                  ), //i
    .io_randW       (randW_x_15_10[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_10_15[14:0]             ), //i
    .io_ofm         (ofm_x_10_16[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_474_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_474_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_474_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_474_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_474_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_474_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_474_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_474_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_474_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_474_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_474_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_474_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_474_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_475 (
    .io_mac_done    (uSystolicPE_475_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_475_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_475_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_475_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_475_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_475_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_475_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_15_11                   ), //i
    .io_ifm_dff     (ifm_dff_x_15_11                    ), //i
    .io_wght_sign   (wght_sign_x_11_15                  ), //i
    .io_randW       (randW_x_15_11[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_11_15[14:0]             ), //i
    .io_ofm         (ofm_x_11_16[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_475_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_475_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_475_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_475_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_475_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_475_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_475_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_475_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_475_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_475_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_475_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_475_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_475_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_476 (
    .io_mac_done    (uSystolicPE_476_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_476_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_476_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_476_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_476_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_476_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_476_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_15_12                   ), //i
    .io_ifm_dff     (ifm_dff_x_15_12                    ), //i
    .io_wght_sign   (wght_sign_x_12_15                  ), //i
    .io_randW       (randW_x_15_12[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_12_15[14:0]             ), //i
    .io_ofm         (ofm_x_12_16[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_476_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_476_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_476_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_476_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_476_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_476_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_476_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_476_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_476_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_476_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_476_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_476_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_476_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_477 (
    .io_mac_done    (uSystolicPE_477_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_477_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_477_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_477_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_477_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_477_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_477_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_15_13                   ), //i
    .io_ifm_dff     (ifm_dff_x_15_13                    ), //i
    .io_wght_sign   (wght_sign_x_13_15                  ), //i
    .io_randW       (randW_x_15_13[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_13_15[14:0]             ), //i
    .io_ofm         (ofm_x_13_16[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_477_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_477_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_477_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_477_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_477_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_477_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_477_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_477_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_477_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_477_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_477_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_477_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_477_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_478 (
    .io_mac_done    (uSystolicPE_478_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_478_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_478_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_478_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_478_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_478_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_478_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_15_14                   ), //i
    .io_ifm_dff     (ifm_dff_x_15_14                    ), //i
    .io_wght_sign   (wght_sign_x_14_15                  ), //i
    .io_randW       (randW_x_15_14[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_14_15[14:0]             ), //i
    .io_ofm         (ofm_x_14_16[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_478_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_478_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_478_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_478_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_478_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_478_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_478_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_478_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_478_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_478_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_478_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_478_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_478_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  uSystolicPE uSystolicPE_479 (
    .io_mac_done    (uSystolicPE_479_io_mac_done        ), //i
    .io_enable_i    (uSystolicPE_479_io_enable_i        ), //i
    .io_clear_i     (uSystolicPE_479_io_clear_i         ), //i
    .io_enable_w    (uSystolicPE_479_io_enable_w        ), //i
    .io_clear_w     (uSystolicPE_479_io_clear_w         ), //i
    .io_enable_o    (uSystolicPE_479_io_enable_o        ), //i
    .io_clear_o     (uSystolicPE_479_io_clear_o         ), //i
    .io_ifm_sign    (ifm_sign_x_15_15                   ), //i
    .io_ifm_dff     (ifm_dff_x_15_15                    ), //i
    .io_wght_sign   (wght_sign_x_15_15                  ), //i
    .io_randW       (randW_x_15_15[14:0]                ), //i
    .io_wght_abs    (wght_abs_x_15_15[14:0]             ), //i
    .io_ofm         (ofm_x_15_16[31:0]                  ), //i
    .io_mac_done_d  (uSystolicPE_479_io_mac_done_d      ), //o
    .io_enable_i_d  (uSystolicPE_479_io_enable_i_d      ), //o
    .io_clear_i_d   (uSystolicPE_479_io_clear_i_d       ), //o
    .io_enable_w_d  (uSystolicPE_479_io_enable_w_d      ), //o
    .io_clear_w_d   (uSystolicPE_479_io_clear_w_d       ), //o
    .io_enable_o_d  (uSystolicPE_479_io_enable_o_d      ), //o
    .io_clear_o_d   (uSystolicPE_479_io_clear_o_d       ), //o
    .io_ifm_sign_d  (uSystolicPE_479_io_ifm_sign_d      ), //o
    .io_ifm_dff_d   (uSystolicPE_479_io_ifm_dff_d       ), //o
    .io_wght_sign_d (uSystolicPE_479_io_wght_sign_d     ), //o
    .io_randW_d     (uSystolicPE_479_io_randW_d[14:0]   ), //o
    .io_wght_abs_d  (uSystolicPE_479_io_wght_abs_d[14:0]), //o
    .io_ofm_d       (uSystolicPE_479_io_ofm_d[31:0]     ), //o
    .clk            (clk                                ), //i
    .reset          (reset                              )  //i
  );
  always @(*) begin
    enable_i_x_0[0] = io_enable_i[0];
    enable_i_x_0[1] = uSystolicPEBorder_16_io_enable_i_d;
    enable_i_x_0[2] = uSystolicPE_240_io_enable_i_d;
    enable_i_x_0[3] = uSystolicPE_241_io_enable_i_d;
    enable_i_x_0[4] = uSystolicPE_242_io_enable_i_d;
    enable_i_x_0[5] = uSystolicPE_243_io_enable_i_d;
    enable_i_x_0[6] = uSystolicPE_244_io_enable_i_d;
    enable_i_x_0[7] = uSystolicPE_245_io_enable_i_d;
    enable_i_x_0[8] = uSystolicPE_246_io_enable_i_d;
    enable_i_x_0[9] = uSystolicPE_247_io_enable_i_d;
    enable_i_x_0[10] = uSystolicPE_248_io_enable_i_d;
    enable_i_x_0[11] = uSystolicPE_249_io_enable_i_d;
    enable_i_x_0[12] = uSystolicPE_250_io_enable_i_d;
    enable_i_x_0[13] = uSystolicPE_251_io_enable_i_d;
    enable_i_x_0[14] = uSystolicPE_252_io_enable_i_d;
    enable_i_x_0[15] = uSystolicPE_253_io_enable_i_d;
    enable_i_x_0[16] = uSystolicPE_254_io_enable_i_d;
  end

  always @(*) begin
    clear_i_x_0[0] = io_clear_i[0];
    clear_i_x_0[1] = uSystolicPEBorder_16_io_clear_i_d;
    clear_i_x_0[2] = uSystolicPE_240_io_clear_i_d;
    clear_i_x_0[3] = uSystolicPE_241_io_clear_i_d;
    clear_i_x_0[4] = uSystolicPE_242_io_clear_i_d;
    clear_i_x_0[5] = uSystolicPE_243_io_clear_i_d;
    clear_i_x_0[6] = uSystolicPE_244_io_clear_i_d;
    clear_i_x_0[7] = uSystolicPE_245_io_clear_i_d;
    clear_i_x_0[8] = uSystolicPE_246_io_clear_i_d;
    clear_i_x_0[9] = uSystolicPE_247_io_clear_i_d;
    clear_i_x_0[10] = uSystolicPE_248_io_clear_i_d;
    clear_i_x_0[11] = uSystolicPE_249_io_clear_i_d;
    clear_i_x_0[12] = uSystolicPE_250_io_clear_i_d;
    clear_i_x_0[13] = uSystolicPE_251_io_clear_i_d;
    clear_i_x_0[14] = uSystolicPE_252_io_clear_i_d;
    clear_i_x_0[15] = uSystolicPE_253_io_clear_i_d;
    clear_i_x_0[16] = uSystolicPE_254_io_clear_i_d;
  end

  always @(*) begin
    mac_done_x_0[0] = io_mac_done[0];
    mac_done_x_0[1] = uSystolicPEBorder_16_io_mac_done_d;
    mac_done_x_0[2] = uSystolicPE_240_io_mac_done_d;
    mac_done_x_0[3] = uSystolicPE_241_io_mac_done_d;
    mac_done_x_0[4] = uSystolicPE_242_io_mac_done_d;
    mac_done_x_0[5] = uSystolicPE_243_io_mac_done_d;
    mac_done_x_0[6] = uSystolicPE_244_io_mac_done_d;
    mac_done_x_0[7] = uSystolicPE_245_io_mac_done_d;
    mac_done_x_0[8] = uSystolicPE_246_io_mac_done_d;
    mac_done_x_0[9] = uSystolicPE_247_io_mac_done_d;
    mac_done_x_0[10] = uSystolicPE_248_io_mac_done_d;
    mac_done_x_0[11] = uSystolicPE_249_io_mac_done_d;
    mac_done_x_0[12] = uSystolicPE_250_io_mac_done_d;
    mac_done_x_0[13] = uSystolicPE_251_io_mac_done_d;
    mac_done_x_0[14] = uSystolicPE_252_io_mac_done_d;
    mac_done_x_0[15] = uSystolicPE_253_io_mac_done_d;
    mac_done_x_0[16] = uSystolicPE_254_io_mac_done_d;
  end

  always @(*) begin
    enable_w_x_0[0] = io_enable_w[0];
    enable_w_x_0[1] = uSystolicPEBorder_16_io_enable_w_d;
    enable_w_x_0[2] = uSystolicPEBorder_17_io_enable_w_d;
    enable_w_x_0[3] = uSystolicPEBorder_18_io_enable_w_d;
    enable_w_x_0[4] = uSystolicPEBorder_19_io_enable_w_d;
    enable_w_x_0[5] = uSystolicPEBorder_20_io_enable_w_d;
    enable_w_x_0[6] = uSystolicPEBorder_21_io_enable_w_d;
    enable_w_x_0[7] = uSystolicPEBorder_22_io_enable_w_d;
    enable_w_x_0[8] = uSystolicPEBorder_23_io_enable_w_d;
    enable_w_x_0[9] = uSystolicPEBorder_24_io_enable_w_d;
    enable_w_x_0[10] = uSystolicPEBorder_25_io_enable_w_d;
    enable_w_x_0[11] = uSystolicPEBorder_26_io_enable_w_d;
    enable_w_x_0[12] = uSystolicPEBorder_27_io_enable_w_d;
    enable_w_x_0[13] = uSystolicPEBorder_28_io_enable_w_d;
    enable_w_x_0[14] = uSystolicPEBorder_29_io_enable_w_d;
    enable_w_x_0[15] = uSystolicPEBorder_30_io_enable_w_d;
    enable_w_x_0[16] = uSystolicPEBorder_31_io_enable_w_d;
  end

  always @(*) begin
    clear_w_x_0[0] = io_clear_w[0];
    clear_w_x_0[1] = uSystolicPEBorder_16_io_clear_w_d;
    clear_w_x_0[2] = uSystolicPEBorder_17_io_clear_w_d;
    clear_w_x_0[3] = uSystolicPEBorder_18_io_clear_w_d;
    clear_w_x_0[4] = uSystolicPEBorder_19_io_clear_w_d;
    clear_w_x_0[5] = uSystolicPEBorder_20_io_clear_w_d;
    clear_w_x_0[6] = uSystolicPEBorder_21_io_clear_w_d;
    clear_w_x_0[7] = uSystolicPEBorder_22_io_clear_w_d;
    clear_w_x_0[8] = uSystolicPEBorder_23_io_clear_w_d;
    clear_w_x_0[9] = uSystolicPEBorder_24_io_clear_w_d;
    clear_w_x_0[10] = uSystolicPEBorder_25_io_clear_w_d;
    clear_w_x_0[11] = uSystolicPEBorder_26_io_clear_w_d;
    clear_w_x_0[12] = uSystolicPEBorder_27_io_clear_w_d;
    clear_w_x_0[13] = uSystolicPEBorder_28_io_clear_w_d;
    clear_w_x_0[14] = uSystolicPEBorder_29_io_clear_w_d;
    clear_w_x_0[15] = uSystolicPEBorder_30_io_clear_w_d;
    clear_w_x_0[16] = uSystolicPEBorder_31_io_clear_w_d;
  end

  assign wght_sign_x_0_0 = io_wght_sign[0];
  assign wght_abs_x_0_0 = io_wght_abs_0;
  always @(*) begin
    enable_o_x_0[16] = io_enable_o[0];
    enable_o_x_0[0] = uSystolicPEBorder_16_io_enable_o_d;
    enable_o_x_0[1] = uSystolicPEBorder_17_io_enable_o_d;
    enable_o_x_0[2] = uSystolicPEBorder_18_io_enable_o_d;
    enable_o_x_0[3] = uSystolicPEBorder_19_io_enable_o_d;
    enable_o_x_0[4] = uSystolicPEBorder_20_io_enable_o_d;
    enable_o_x_0[5] = uSystolicPEBorder_21_io_enable_o_d;
    enable_o_x_0[6] = uSystolicPEBorder_22_io_enable_o_d;
    enable_o_x_0[7] = uSystolicPEBorder_23_io_enable_o_d;
    enable_o_x_0[8] = uSystolicPEBorder_24_io_enable_o_d;
    enable_o_x_0[9] = uSystolicPEBorder_25_io_enable_o_d;
    enable_o_x_0[10] = uSystolicPEBorder_26_io_enable_o_d;
    enable_o_x_0[11] = uSystolicPEBorder_27_io_enable_o_d;
    enable_o_x_0[12] = uSystolicPEBorder_28_io_enable_o_d;
    enable_o_x_0[13] = uSystolicPEBorder_29_io_enable_o_d;
    enable_o_x_0[14] = uSystolicPEBorder_30_io_enable_o_d;
    enable_o_x_0[15] = uSystolicPEBorder_31_io_enable_o_d;
  end

  always @(*) begin
    clear_o_x_0[16] = io_clear_o[0];
    clear_o_x_0[0] = uSystolicPEBorder_16_io_clear_o_d;
    clear_o_x_0[1] = uSystolicPEBorder_17_io_clear_o_d;
    clear_o_x_0[2] = uSystolicPEBorder_18_io_clear_o_d;
    clear_o_x_0[3] = uSystolicPEBorder_19_io_clear_o_d;
    clear_o_x_0[4] = uSystolicPEBorder_20_io_clear_o_d;
    clear_o_x_0[5] = uSystolicPEBorder_21_io_clear_o_d;
    clear_o_x_0[6] = uSystolicPEBorder_22_io_clear_o_d;
    clear_o_x_0[7] = uSystolicPEBorder_23_io_clear_o_d;
    clear_o_x_0[8] = uSystolicPEBorder_24_io_clear_o_d;
    clear_o_x_0[9] = uSystolicPEBorder_25_io_clear_o_d;
    clear_o_x_0[10] = uSystolicPEBorder_26_io_clear_o_d;
    clear_o_x_0[11] = uSystolicPEBorder_27_io_clear_o_d;
    clear_o_x_0[12] = uSystolicPEBorder_28_io_clear_o_d;
    clear_o_x_0[13] = uSystolicPEBorder_29_io_clear_o_d;
    clear_o_x_0[14] = uSystolicPEBorder_30_io_clear_o_d;
    clear_o_x_0[15] = uSystolicPEBorder_31_io_clear_o_d;
  end

  assign io_ofm_0 = ofm_x_0_0;
  assign ofm_x_0_16 = 32'h00000000;
  always @(*) begin
    enable_i_x_1[0] = io_enable_i[1];
    enable_i_x_1[1] = uSystolicPEBorder_17_io_enable_i_d;
    enable_i_x_1[2] = uSystolicPE_255_io_enable_i_d;
    enable_i_x_1[3] = uSystolicPE_256_io_enable_i_d;
    enable_i_x_1[4] = uSystolicPE_257_io_enable_i_d;
    enable_i_x_1[5] = uSystolicPE_258_io_enable_i_d;
    enable_i_x_1[6] = uSystolicPE_259_io_enable_i_d;
    enable_i_x_1[7] = uSystolicPE_260_io_enable_i_d;
    enable_i_x_1[8] = uSystolicPE_261_io_enable_i_d;
    enable_i_x_1[9] = uSystolicPE_262_io_enable_i_d;
    enable_i_x_1[10] = uSystolicPE_263_io_enable_i_d;
    enable_i_x_1[11] = uSystolicPE_264_io_enable_i_d;
    enable_i_x_1[12] = uSystolicPE_265_io_enable_i_d;
    enable_i_x_1[13] = uSystolicPE_266_io_enable_i_d;
    enable_i_x_1[14] = uSystolicPE_267_io_enable_i_d;
    enable_i_x_1[15] = uSystolicPE_268_io_enable_i_d;
    enable_i_x_1[16] = uSystolicPE_269_io_enable_i_d;
  end

  always @(*) begin
    clear_i_x_1[0] = io_clear_i[1];
    clear_i_x_1[1] = uSystolicPEBorder_17_io_clear_i_d;
    clear_i_x_1[2] = uSystolicPE_255_io_clear_i_d;
    clear_i_x_1[3] = uSystolicPE_256_io_clear_i_d;
    clear_i_x_1[4] = uSystolicPE_257_io_clear_i_d;
    clear_i_x_1[5] = uSystolicPE_258_io_clear_i_d;
    clear_i_x_1[6] = uSystolicPE_259_io_clear_i_d;
    clear_i_x_1[7] = uSystolicPE_260_io_clear_i_d;
    clear_i_x_1[8] = uSystolicPE_261_io_clear_i_d;
    clear_i_x_1[9] = uSystolicPE_262_io_clear_i_d;
    clear_i_x_1[10] = uSystolicPE_263_io_clear_i_d;
    clear_i_x_1[11] = uSystolicPE_264_io_clear_i_d;
    clear_i_x_1[12] = uSystolicPE_265_io_clear_i_d;
    clear_i_x_1[13] = uSystolicPE_266_io_clear_i_d;
    clear_i_x_1[14] = uSystolicPE_267_io_clear_i_d;
    clear_i_x_1[15] = uSystolicPE_268_io_clear_i_d;
    clear_i_x_1[16] = uSystolicPE_269_io_clear_i_d;
  end

  always @(*) begin
    mac_done_x_1[0] = io_mac_done[1];
    mac_done_x_1[1] = uSystolicPEBorder_17_io_mac_done_d;
    mac_done_x_1[2] = uSystolicPE_255_io_mac_done_d;
    mac_done_x_1[3] = uSystolicPE_256_io_mac_done_d;
    mac_done_x_1[4] = uSystolicPE_257_io_mac_done_d;
    mac_done_x_1[5] = uSystolicPE_258_io_mac_done_d;
    mac_done_x_1[6] = uSystolicPE_259_io_mac_done_d;
    mac_done_x_1[7] = uSystolicPE_260_io_mac_done_d;
    mac_done_x_1[8] = uSystolicPE_261_io_mac_done_d;
    mac_done_x_1[9] = uSystolicPE_262_io_mac_done_d;
    mac_done_x_1[10] = uSystolicPE_263_io_mac_done_d;
    mac_done_x_1[11] = uSystolicPE_264_io_mac_done_d;
    mac_done_x_1[12] = uSystolicPE_265_io_mac_done_d;
    mac_done_x_1[13] = uSystolicPE_266_io_mac_done_d;
    mac_done_x_1[14] = uSystolicPE_267_io_mac_done_d;
    mac_done_x_1[15] = uSystolicPE_268_io_mac_done_d;
    mac_done_x_1[16] = uSystolicPE_269_io_mac_done_d;
  end

  always @(*) begin
    enable_w_x_1[0] = io_enable_w[1];
    enable_w_x_1[1] = uSystolicPE_240_io_enable_w_d;
    enable_w_x_1[2] = uSystolicPE_255_io_enable_w_d;
    enable_w_x_1[3] = uSystolicPE_270_io_enable_w_d;
    enable_w_x_1[4] = uSystolicPE_285_io_enable_w_d;
    enable_w_x_1[5] = uSystolicPE_300_io_enable_w_d;
    enable_w_x_1[6] = uSystolicPE_315_io_enable_w_d;
    enable_w_x_1[7] = uSystolicPE_330_io_enable_w_d;
    enable_w_x_1[8] = uSystolicPE_345_io_enable_w_d;
    enable_w_x_1[9] = uSystolicPE_360_io_enable_w_d;
    enable_w_x_1[10] = uSystolicPE_375_io_enable_w_d;
    enable_w_x_1[11] = uSystolicPE_390_io_enable_w_d;
    enable_w_x_1[12] = uSystolicPE_405_io_enable_w_d;
    enable_w_x_1[13] = uSystolicPE_420_io_enable_w_d;
    enable_w_x_1[14] = uSystolicPE_435_io_enable_w_d;
    enable_w_x_1[15] = uSystolicPE_450_io_enable_w_d;
    enable_w_x_1[16] = uSystolicPE_465_io_enable_w_d;
  end

  always @(*) begin
    clear_w_x_1[0] = io_clear_w[1];
    clear_w_x_1[1] = uSystolicPE_240_io_clear_w_d;
    clear_w_x_1[2] = uSystolicPE_255_io_clear_w_d;
    clear_w_x_1[3] = uSystolicPE_270_io_clear_w_d;
    clear_w_x_1[4] = uSystolicPE_285_io_clear_w_d;
    clear_w_x_1[5] = uSystolicPE_300_io_clear_w_d;
    clear_w_x_1[6] = uSystolicPE_315_io_clear_w_d;
    clear_w_x_1[7] = uSystolicPE_330_io_clear_w_d;
    clear_w_x_1[8] = uSystolicPE_345_io_clear_w_d;
    clear_w_x_1[9] = uSystolicPE_360_io_clear_w_d;
    clear_w_x_1[10] = uSystolicPE_375_io_clear_w_d;
    clear_w_x_1[11] = uSystolicPE_390_io_clear_w_d;
    clear_w_x_1[12] = uSystolicPE_405_io_clear_w_d;
    clear_w_x_1[13] = uSystolicPE_420_io_clear_w_d;
    clear_w_x_1[14] = uSystolicPE_435_io_clear_w_d;
    clear_w_x_1[15] = uSystolicPE_450_io_clear_w_d;
    clear_w_x_1[16] = uSystolicPE_465_io_clear_w_d;
  end

  assign wght_sign_x_1_0 = io_wght_sign[1];
  assign wght_abs_x_1_0 = io_wght_abs_1;
  always @(*) begin
    enable_o_x_1[16] = io_enable_o[1];
    enable_o_x_1[0] = uSystolicPE_240_io_enable_o_d;
    enable_o_x_1[1] = uSystolicPE_255_io_enable_o_d;
    enable_o_x_1[2] = uSystolicPE_270_io_enable_o_d;
    enable_o_x_1[3] = uSystolicPE_285_io_enable_o_d;
    enable_o_x_1[4] = uSystolicPE_300_io_enable_o_d;
    enable_o_x_1[5] = uSystolicPE_315_io_enable_o_d;
    enable_o_x_1[6] = uSystolicPE_330_io_enable_o_d;
    enable_o_x_1[7] = uSystolicPE_345_io_enable_o_d;
    enable_o_x_1[8] = uSystolicPE_360_io_enable_o_d;
    enable_o_x_1[9] = uSystolicPE_375_io_enable_o_d;
    enable_o_x_1[10] = uSystolicPE_390_io_enable_o_d;
    enable_o_x_1[11] = uSystolicPE_405_io_enable_o_d;
    enable_o_x_1[12] = uSystolicPE_420_io_enable_o_d;
    enable_o_x_1[13] = uSystolicPE_435_io_enable_o_d;
    enable_o_x_1[14] = uSystolicPE_450_io_enable_o_d;
    enable_o_x_1[15] = uSystolicPE_465_io_enable_o_d;
  end

  always @(*) begin
    clear_o_x_1[16] = io_clear_o[1];
    clear_o_x_1[0] = uSystolicPE_240_io_clear_o_d;
    clear_o_x_1[1] = uSystolicPE_255_io_clear_o_d;
    clear_o_x_1[2] = uSystolicPE_270_io_clear_o_d;
    clear_o_x_1[3] = uSystolicPE_285_io_clear_o_d;
    clear_o_x_1[4] = uSystolicPE_300_io_clear_o_d;
    clear_o_x_1[5] = uSystolicPE_315_io_clear_o_d;
    clear_o_x_1[6] = uSystolicPE_330_io_clear_o_d;
    clear_o_x_1[7] = uSystolicPE_345_io_clear_o_d;
    clear_o_x_1[8] = uSystolicPE_360_io_clear_o_d;
    clear_o_x_1[9] = uSystolicPE_375_io_clear_o_d;
    clear_o_x_1[10] = uSystolicPE_390_io_clear_o_d;
    clear_o_x_1[11] = uSystolicPE_405_io_clear_o_d;
    clear_o_x_1[12] = uSystolicPE_420_io_clear_o_d;
    clear_o_x_1[13] = uSystolicPE_435_io_clear_o_d;
    clear_o_x_1[14] = uSystolicPE_450_io_clear_o_d;
    clear_o_x_1[15] = uSystolicPE_465_io_clear_o_d;
  end

  assign io_ofm_1 = ofm_x_1_0;
  assign ofm_x_1_16 = 32'h00000000;
  always @(*) begin
    enable_i_x_2[0] = io_enable_i[2];
    enable_i_x_2[1] = uSystolicPEBorder_18_io_enable_i_d;
    enable_i_x_2[2] = uSystolicPE_270_io_enable_i_d;
    enable_i_x_2[3] = uSystolicPE_271_io_enable_i_d;
    enable_i_x_2[4] = uSystolicPE_272_io_enable_i_d;
    enable_i_x_2[5] = uSystolicPE_273_io_enable_i_d;
    enable_i_x_2[6] = uSystolicPE_274_io_enable_i_d;
    enable_i_x_2[7] = uSystolicPE_275_io_enable_i_d;
    enable_i_x_2[8] = uSystolicPE_276_io_enable_i_d;
    enable_i_x_2[9] = uSystolicPE_277_io_enable_i_d;
    enable_i_x_2[10] = uSystolicPE_278_io_enable_i_d;
    enable_i_x_2[11] = uSystolicPE_279_io_enable_i_d;
    enable_i_x_2[12] = uSystolicPE_280_io_enable_i_d;
    enable_i_x_2[13] = uSystolicPE_281_io_enable_i_d;
    enable_i_x_2[14] = uSystolicPE_282_io_enable_i_d;
    enable_i_x_2[15] = uSystolicPE_283_io_enable_i_d;
    enable_i_x_2[16] = uSystolicPE_284_io_enable_i_d;
  end

  always @(*) begin
    clear_i_x_2[0] = io_clear_i[2];
    clear_i_x_2[1] = uSystolicPEBorder_18_io_clear_i_d;
    clear_i_x_2[2] = uSystolicPE_270_io_clear_i_d;
    clear_i_x_2[3] = uSystolicPE_271_io_clear_i_d;
    clear_i_x_2[4] = uSystolicPE_272_io_clear_i_d;
    clear_i_x_2[5] = uSystolicPE_273_io_clear_i_d;
    clear_i_x_2[6] = uSystolicPE_274_io_clear_i_d;
    clear_i_x_2[7] = uSystolicPE_275_io_clear_i_d;
    clear_i_x_2[8] = uSystolicPE_276_io_clear_i_d;
    clear_i_x_2[9] = uSystolicPE_277_io_clear_i_d;
    clear_i_x_2[10] = uSystolicPE_278_io_clear_i_d;
    clear_i_x_2[11] = uSystolicPE_279_io_clear_i_d;
    clear_i_x_2[12] = uSystolicPE_280_io_clear_i_d;
    clear_i_x_2[13] = uSystolicPE_281_io_clear_i_d;
    clear_i_x_2[14] = uSystolicPE_282_io_clear_i_d;
    clear_i_x_2[15] = uSystolicPE_283_io_clear_i_d;
    clear_i_x_2[16] = uSystolicPE_284_io_clear_i_d;
  end

  always @(*) begin
    mac_done_x_2[0] = io_mac_done[2];
    mac_done_x_2[1] = uSystolicPEBorder_18_io_mac_done_d;
    mac_done_x_2[2] = uSystolicPE_270_io_mac_done_d;
    mac_done_x_2[3] = uSystolicPE_271_io_mac_done_d;
    mac_done_x_2[4] = uSystolicPE_272_io_mac_done_d;
    mac_done_x_2[5] = uSystolicPE_273_io_mac_done_d;
    mac_done_x_2[6] = uSystolicPE_274_io_mac_done_d;
    mac_done_x_2[7] = uSystolicPE_275_io_mac_done_d;
    mac_done_x_2[8] = uSystolicPE_276_io_mac_done_d;
    mac_done_x_2[9] = uSystolicPE_277_io_mac_done_d;
    mac_done_x_2[10] = uSystolicPE_278_io_mac_done_d;
    mac_done_x_2[11] = uSystolicPE_279_io_mac_done_d;
    mac_done_x_2[12] = uSystolicPE_280_io_mac_done_d;
    mac_done_x_2[13] = uSystolicPE_281_io_mac_done_d;
    mac_done_x_2[14] = uSystolicPE_282_io_mac_done_d;
    mac_done_x_2[15] = uSystolicPE_283_io_mac_done_d;
    mac_done_x_2[16] = uSystolicPE_284_io_mac_done_d;
  end

  always @(*) begin
    enable_w_x_2[0] = io_enable_w[2];
    enable_w_x_2[1] = uSystolicPE_241_io_enable_w_d;
    enable_w_x_2[2] = uSystolicPE_256_io_enable_w_d;
    enable_w_x_2[3] = uSystolicPE_271_io_enable_w_d;
    enable_w_x_2[4] = uSystolicPE_286_io_enable_w_d;
    enable_w_x_2[5] = uSystolicPE_301_io_enable_w_d;
    enable_w_x_2[6] = uSystolicPE_316_io_enable_w_d;
    enable_w_x_2[7] = uSystolicPE_331_io_enable_w_d;
    enable_w_x_2[8] = uSystolicPE_346_io_enable_w_d;
    enable_w_x_2[9] = uSystolicPE_361_io_enable_w_d;
    enable_w_x_2[10] = uSystolicPE_376_io_enable_w_d;
    enable_w_x_2[11] = uSystolicPE_391_io_enable_w_d;
    enable_w_x_2[12] = uSystolicPE_406_io_enable_w_d;
    enable_w_x_2[13] = uSystolicPE_421_io_enable_w_d;
    enable_w_x_2[14] = uSystolicPE_436_io_enable_w_d;
    enable_w_x_2[15] = uSystolicPE_451_io_enable_w_d;
    enable_w_x_2[16] = uSystolicPE_466_io_enable_w_d;
  end

  always @(*) begin
    clear_w_x_2[0] = io_clear_w[2];
    clear_w_x_2[1] = uSystolicPE_241_io_clear_w_d;
    clear_w_x_2[2] = uSystolicPE_256_io_clear_w_d;
    clear_w_x_2[3] = uSystolicPE_271_io_clear_w_d;
    clear_w_x_2[4] = uSystolicPE_286_io_clear_w_d;
    clear_w_x_2[5] = uSystolicPE_301_io_clear_w_d;
    clear_w_x_2[6] = uSystolicPE_316_io_clear_w_d;
    clear_w_x_2[7] = uSystolicPE_331_io_clear_w_d;
    clear_w_x_2[8] = uSystolicPE_346_io_clear_w_d;
    clear_w_x_2[9] = uSystolicPE_361_io_clear_w_d;
    clear_w_x_2[10] = uSystolicPE_376_io_clear_w_d;
    clear_w_x_2[11] = uSystolicPE_391_io_clear_w_d;
    clear_w_x_2[12] = uSystolicPE_406_io_clear_w_d;
    clear_w_x_2[13] = uSystolicPE_421_io_clear_w_d;
    clear_w_x_2[14] = uSystolicPE_436_io_clear_w_d;
    clear_w_x_2[15] = uSystolicPE_451_io_clear_w_d;
    clear_w_x_2[16] = uSystolicPE_466_io_clear_w_d;
  end

  assign wght_sign_x_2_0 = io_wght_sign[2];
  assign wght_abs_x_2_0 = io_wght_abs_2;
  always @(*) begin
    enable_o_x_2[16] = io_enable_o[2];
    enable_o_x_2[0] = uSystolicPE_241_io_enable_o_d;
    enable_o_x_2[1] = uSystolicPE_256_io_enable_o_d;
    enable_o_x_2[2] = uSystolicPE_271_io_enable_o_d;
    enable_o_x_2[3] = uSystolicPE_286_io_enable_o_d;
    enable_o_x_2[4] = uSystolicPE_301_io_enable_o_d;
    enable_o_x_2[5] = uSystolicPE_316_io_enable_o_d;
    enable_o_x_2[6] = uSystolicPE_331_io_enable_o_d;
    enable_o_x_2[7] = uSystolicPE_346_io_enable_o_d;
    enable_o_x_2[8] = uSystolicPE_361_io_enable_o_d;
    enable_o_x_2[9] = uSystolicPE_376_io_enable_o_d;
    enable_o_x_2[10] = uSystolicPE_391_io_enable_o_d;
    enable_o_x_2[11] = uSystolicPE_406_io_enable_o_d;
    enable_o_x_2[12] = uSystolicPE_421_io_enable_o_d;
    enable_o_x_2[13] = uSystolicPE_436_io_enable_o_d;
    enable_o_x_2[14] = uSystolicPE_451_io_enable_o_d;
    enable_o_x_2[15] = uSystolicPE_466_io_enable_o_d;
  end

  always @(*) begin
    clear_o_x_2[16] = io_clear_o[2];
    clear_o_x_2[0] = uSystolicPE_241_io_clear_o_d;
    clear_o_x_2[1] = uSystolicPE_256_io_clear_o_d;
    clear_o_x_2[2] = uSystolicPE_271_io_clear_o_d;
    clear_o_x_2[3] = uSystolicPE_286_io_clear_o_d;
    clear_o_x_2[4] = uSystolicPE_301_io_clear_o_d;
    clear_o_x_2[5] = uSystolicPE_316_io_clear_o_d;
    clear_o_x_2[6] = uSystolicPE_331_io_clear_o_d;
    clear_o_x_2[7] = uSystolicPE_346_io_clear_o_d;
    clear_o_x_2[8] = uSystolicPE_361_io_clear_o_d;
    clear_o_x_2[9] = uSystolicPE_376_io_clear_o_d;
    clear_o_x_2[10] = uSystolicPE_391_io_clear_o_d;
    clear_o_x_2[11] = uSystolicPE_406_io_clear_o_d;
    clear_o_x_2[12] = uSystolicPE_421_io_clear_o_d;
    clear_o_x_2[13] = uSystolicPE_436_io_clear_o_d;
    clear_o_x_2[14] = uSystolicPE_451_io_clear_o_d;
    clear_o_x_2[15] = uSystolicPE_466_io_clear_o_d;
  end

  assign io_ofm_2 = ofm_x_2_0;
  assign ofm_x_2_16 = 32'h00000000;
  always @(*) begin
    enable_i_x_3[0] = io_enable_i[3];
    enable_i_x_3[1] = uSystolicPEBorder_19_io_enable_i_d;
    enable_i_x_3[2] = uSystolicPE_285_io_enable_i_d;
    enable_i_x_3[3] = uSystolicPE_286_io_enable_i_d;
    enable_i_x_3[4] = uSystolicPE_287_io_enable_i_d;
    enable_i_x_3[5] = uSystolicPE_288_io_enable_i_d;
    enable_i_x_3[6] = uSystolicPE_289_io_enable_i_d;
    enable_i_x_3[7] = uSystolicPE_290_io_enable_i_d;
    enable_i_x_3[8] = uSystolicPE_291_io_enable_i_d;
    enable_i_x_3[9] = uSystolicPE_292_io_enable_i_d;
    enable_i_x_3[10] = uSystolicPE_293_io_enable_i_d;
    enable_i_x_3[11] = uSystolicPE_294_io_enable_i_d;
    enable_i_x_3[12] = uSystolicPE_295_io_enable_i_d;
    enable_i_x_3[13] = uSystolicPE_296_io_enable_i_d;
    enable_i_x_3[14] = uSystolicPE_297_io_enable_i_d;
    enable_i_x_3[15] = uSystolicPE_298_io_enable_i_d;
    enable_i_x_3[16] = uSystolicPE_299_io_enable_i_d;
  end

  always @(*) begin
    clear_i_x_3[0] = io_clear_i[3];
    clear_i_x_3[1] = uSystolicPEBorder_19_io_clear_i_d;
    clear_i_x_3[2] = uSystolicPE_285_io_clear_i_d;
    clear_i_x_3[3] = uSystolicPE_286_io_clear_i_d;
    clear_i_x_3[4] = uSystolicPE_287_io_clear_i_d;
    clear_i_x_3[5] = uSystolicPE_288_io_clear_i_d;
    clear_i_x_3[6] = uSystolicPE_289_io_clear_i_d;
    clear_i_x_3[7] = uSystolicPE_290_io_clear_i_d;
    clear_i_x_3[8] = uSystolicPE_291_io_clear_i_d;
    clear_i_x_3[9] = uSystolicPE_292_io_clear_i_d;
    clear_i_x_3[10] = uSystolicPE_293_io_clear_i_d;
    clear_i_x_3[11] = uSystolicPE_294_io_clear_i_d;
    clear_i_x_3[12] = uSystolicPE_295_io_clear_i_d;
    clear_i_x_3[13] = uSystolicPE_296_io_clear_i_d;
    clear_i_x_3[14] = uSystolicPE_297_io_clear_i_d;
    clear_i_x_3[15] = uSystolicPE_298_io_clear_i_d;
    clear_i_x_3[16] = uSystolicPE_299_io_clear_i_d;
  end

  always @(*) begin
    mac_done_x_3[0] = io_mac_done[3];
    mac_done_x_3[1] = uSystolicPEBorder_19_io_mac_done_d;
    mac_done_x_3[2] = uSystolicPE_285_io_mac_done_d;
    mac_done_x_3[3] = uSystolicPE_286_io_mac_done_d;
    mac_done_x_3[4] = uSystolicPE_287_io_mac_done_d;
    mac_done_x_3[5] = uSystolicPE_288_io_mac_done_d;
    mac_done_x_3[6] = uSystolicPE_289_io_mac_done_d;
    mac_done_x_3[7] = uSystolicPE_290_io_mac_done_d;
    mac_done_x_3[8] = uSystolicPE_291_io_mac_done_d;
    mac_done_x_3[9] = uSystolicPE_292_io_mac_done_d;
    mac_done_x_3[10] = uSystolicPE_293_io_mac_done_d;
    mac_done_x_3[11] = uSystolicPE_294_io_mac_done_d;
    mac_done_x_3[12] = uSystolicPE_295_io_mac_done_d;
    mac_done_x_3[13] = uSystolicPE_296_io_mac_done_d;
    mac_done_x_3[14] = uSystolicPE_297_io_mac_done_d;
    mac_done_x_3[15] = uSystolicPE_298_io_mac_done_d;
    mac_done_x_3[16] = uSystolicPE_299_io_mac_done_d;
  end

  always @(*) begin
    enable_w_x_3[0] = io_enable_w[3];
    enable_w_x_3[1] = uSystolicPE_242_io_enable_w_d;
    enable_w_x_3[2] = uSystolicPE_257_io_enable_w_d;
    enable_w_x_3[3] = uSystolicPE_272_io_enable_w_d;
    enable_w_x_3[4] = uSystolicPE_287_io_enable_w_d;
    enable_w_x_3[5] = uSystolicPE_302_io_enable_w_d;
    enable_w_x_3[6] = uSystolicPE_317_io_enable_w_d;
    enable_w_x_3[7] = uSystolicPE_332_io_enable_w_d;
    enable_w_x_3[8] = uSystolicPE_347_io_enable_w_d;
    enable_w_x_3[9] = uSystolicPE_362_io_enable_w_d;
    enable_w_x_3[10] = uSystolicPE_377_io_enable_w_d;
    enable_w_x_3[11] = uSystolicPE_392_io_enable_w_d;
    enable_w_x_3[12] = uSystolicPE_407_io_enable_w_d;
    enable_w_x_3[13] = uSystolicPE_422_io_enable_w_d;
    enable_w_x_3[14] = uSystolicPE_437_io_enable_w_d;
    enable_w_x_3[15] = uSystolicPE_452_io_enable_w_d;
    enable_w_x_3[16] = uSystolicPE_467_io_enable_w_d;
  end

  always @(*) begin
    clear_w_x_3[0] = io_clear_w[3];
    clear_w_x_3[1] = uSystolicPE_242_io_clear_w_d;
    clear_w_x_3[2] = uSystolicPE_257_io_clear_w_d;
    clear_w_x_3[3] = uSystolicPE_272_io_clear_w_d;
    clear_w_x_3[4] = uSystolicPE_287_io_clear_w_d;
    clear_w_x_3[5] = uSystolicPE_302_io_clear_w_d;
    clear_w_x_3[6] = uSystolicPE_317_io_clear_w_d;
    clear_w_x_3[7] = uSystolicPE_332_io_clear_w_d;
    clear_w_x_3[8] = uSystolicPE_347_io_clear_w_d;
    clear_w_x_3[9] = uSystolicPE_362_io_clear_w_d;
    clear_w_x_3[10] = uSystolicPE_377_io_clear_w_d;
    clear_w_x_3[11] = uSystolicPE_392_io_clear_w_d;
    clear_w_x_3[12] = uSystolicPE_407_io_clear_w_d;
    clear_w_x_3[13] = uSystolicPE_422_io_clear_w_d;
    clear_w_x_3[14] = uSystolicPE_437_io_clear_w_d;
    clear_w_x_3[15] = uSystolicPE_452_io_clear_w_d;
    clear_w_x_3[16] = uSystolicPE_467_io_clear_w_d;
  end

  assign wght_sign_x_3_0 = io_wght_sign[3];
  assign wght_abs_x_3_0 = io_wght_abs_3;
  always @(*) begin
    enable_o_x_3[16] = io_enable_o[3];
    enable_o_x_3[0] = uSystolicPE_242_io_enable_o_d;
    enable_o_x_3[1] = uSystolicPE_257_io_enable_o_d;
    enable_o_x_3[2] = uSystolicPE_272_io_enable_o_d;
    enable_o_x_3[3] = uSystolicPE_287_io_enable_o_d;
    enable_o_x_3[4] = uSystolicPE_302_io_enable_o_d;
    enable_o_x_3[5] = uSystolicPE_317_io_enable_o_d;
    enable_o_x_3[6] = uSystolicPE_332_io_enable_o_d;
    enable_o_x_3[7] = uSystolicPE_347_io_enable_o_d;
    enable_o_x_3[8] = uSystolicPE_362_io_enable_o_d;
    enable_o_x_3[9] = uSystolicPE_377_io_enable_o_d;
    enable_o_x_3[10] = uSystolicPE_392_io_enable_o_d;
    enable_o_x_3[11] = uSystolicPE_407_io_enable_o_d;
    enable_o_x_3[12] = uSystolicPE_422_io_enable_o_d;
    enable_o_x_3[13] = uSystolicPE_437_io_enable_o_d;
    enable_o_x_3[14] = uSystolicPE_452_io_enable_o_d;
    enable_o_x_3[15] = uSystolicPE_467_io_enable_o_d;
  end

  always @(*) begin
    clear_o_x_3[16] = io_clear_o[3];
    clear_o_x_3[0] = uSystolicPE_242_io_clear_o_d;
    clear_o_x_3[1] = uSystolicPE_257_io_clear_o_d;
    clear_o_x_3[2] = uSystolicPE_272_io_clear_o_d;
    clear_o_x_3[3] = uSystolicPE_287_io_clear_o_d;
    clear_o_x_3[4] = uSystolicPE_302_io_clear_o_d;
    clear_o_x_3[5] = uSystolicPE_317_io_clear_o_d;
    clear_o_x_3[6] = uSystolicPE_332_io_clear_o_d;
    clear_o_x_3[7] = uSystolicPE_347_io_clear_o_d;
    clear_o_x_3[8] = uSystolicPE_362_io_clear_o_d;
    clear_o_x_3[9] = uSystolicPE_377_io_clear_o_d;
    clear_o_x_3[10] = uSystolicPE_392_io_clear_o_d;
    clear_o_x_3[11] = uSystolicPE_407_io_clear_o_d;
    clear_o_x_3[12] = uSystolicPE_422_io_clear_o_d;
    clear_o_x_3[13] = uSystolicPE_437_io_clear_o_d;
    clear_o_x_3[14] = uSystolicPE_452_io_clear_o_d;
    clear_o_x_3[15] = uSystolicPE_467_io_clear_o_d;
  end

  assign io_ofm_3 = ofm_x_3_0;
  assign ofm_x_3_16 = 32'h00000000;
  always @(*) begin
    enable_i_x_4[0] = io_enable_i[4];
    enable_i_x_4[1] = uSystolicPEBorder_20_io_enable_i_d;
    enable_i_x_4[2] = uSystolicPE_300_io_enable_i_d;
    enable_i_x_4[3] = uSystolicPE_301_io_enable_i_d;
    enable_i_x_4[4] = uSystolicPE_302_io_enable_i_d;
    enable_i_x_4[5] = uSystolicPE_303_io_enable_i_d;
    enable_i_x_4[6] = uSystolicPE_304_io_enable_i_d;
    enable_i_x_4[7] = uSystolicPE_305_io_enable_i_d;
    enable_i_x_4[8] = uSystolicPE_306_io_enable_i_d;
    enable_i_x_4[9] = uSystolicPE_307_io_enable_i_d;
    enable_i_x_4[10] = uSystolicPE_308_io_enable_i_d;
    enable_i_x_4[11] = uSystolicPE_309_io_enable_i_d;
    enable_i_x_4[12] = uSystolicPE_310_io_enable_i_d;
    enable_i_x_4[13] = uSystolicPE_311_io_enable_i_d;
    enable_i_x_4[14] = uSystolicPE_312_io_enable_i_d;
    enable_i_x_4[15] = uSystolicPE_313_io_enable_i_d;
    enable_i_x_4[16] = uSystolicPE_314_io_enable_i_d;
  end

  always @(*) begin
    clear_i_x_4[0] = io_clear_i[4];
    clear_i_x_4[1] = uSystolicPEBorder_20_io_clear_i_d;
    clear_i_x_4[2] = uSystolicPE_300_io_clear_i_d;
    clear_i_x_4[3] = uSystolicPE_301_io_clear_i_d;
    clear_i_x_4[4] = uSystolicPE_302_io_clear_i_d;
    clear_i_x_4[5] = uSystolicPE_303_io_clear_i_d;
    clear_i_x_4[6] = uSystolicPE_304_io_clear_i_d;
    clear_i_x_4[7] = uSystolicPE_305_io_clear_i_d;
    clear_i_x_4[8] = uSystolicPE_306_io_clear_i_d;
    clear_i_x_4[9] = uSystolicPE_307_io_clear_i_d;
    clear_i_x_4[10] = uSystolicPE_308_io_clear_i_d;
    clear_i_x_4[11] = uSystolicPE_309_io_clear_i_d;
    clear_i_x_4[12] = uSystolicPE_310_io_clear_i_d;
    clear_i_x_4[13] = uSystolicPE_311_io_clear_i_d;
    clear_i_x_4[14] = uSystolicPE_312_io_clear_i_d;
    clear_i_x_4[15] = uSystolicPE_313_io_clear_i_d;
    clear_i_x_4[16] = uSystolicPE_314_io_clear_i_d;
  end

  always @(*) begin
    mac_done_x_4[0] = io_mac_done[4];
    mac_done_x_4[1] = uSystolicPEBorder_20_io_mac_done_d;
    mac_done_x_4[2] = uSystolicPE_300_io_mac_done_d;
    mac_done_x_4[3] = uSystolicPE_301_io_mac_done_d;
    mac_done_x_4[4] = uSystolicPE_302_io_mac_done_d;
    mac_done_x_4[5] = uSystolicPE_303_io_mac_done_d;
    mac_done_x_4[6] = uSystolicPE_304_io_mac_done_d;
    mac_done_x_4[7] = uSystolicPE_305_io_mac_done_d;
    mac_done_x_4[8] = uSystolicPE_306_io_mac_done_d;
    mac_done_x_4[9] = uSystolicPE_307_io_mac_done_d;
    mac_done_x_4[10] = uSystolicPE_308_io_mac_done_d;
    mac_done_x_4[11] = uSystolicPE_309_io_mac_done_d;
    mac_done_x_4[12] = uSystolicPE_310_io_mac_done_d;
    mac_done_x_4[13] = uSystolicPE_311_io_mac_done_d;
    mac_done_x_4[14] = uSystolicPE_312_io_mac_done_d;
    mac_done_x_4[15] = uSystolicPE_313_io_mac_done_d;
    mac_done_x_4[16] = uSystolicPE_314_io_mac_done_d;
  end

  always @(*) begin
    enable_w_x_4[0] = io_enable_w[4];
    enable_w_x_4[1] = uSystolicPE_243_io_enable_w_d;
    enable_w_x_4[2] = uSystolicPE_258_io_enable_w_d;
    enable_w_x_4[3] = uSystolicPE_273_io_enable_w_d;
    enable_w_x_4[4] = uSystolicPE_288_io_enable_w_d;
    enable_w_x_4[5] = uSystolicPE_303_io_enable_w_d;
    enable_w_x_4[6] = uSystolicPE_318_io_enable_w_d;
    enable_w_x_4[7] = uSystolicPE_333_io_enable_w_d;
    enable_w_x_4[8] = uSystolicPE_348_io_enable_w_d;
    enable_w_x_4[9] = uSystolicPE_363_io_enable_w_d;
    enable_w_x_4[10] = uSystolicPE_378_io_enable_w_d;
    enable_w_x_4[11] = uSystolicPE_393_io_enable_w_d;
    enable_w_x_4[12] = uSystolicPE_408_io_enable_w_d;
    enable_w_x_4[13] = uSystolicPE_423_io_enable_w_d;
    enable_w_x_4[14] = uSystolicPE_438_io_enable_w_d;
    enable_w_x_4[15] = uSystolicPE_453_io_enable_w_d;
    enable_w_x_4[16] = uSystolicPE_468_io_enable_w_d;
  end

  always @(*) begin
    clear_w_x_4[0] = io_clear_w[4];
    clear_w_x_4[1] = uSystolicPE_243_io_clear_w_d;
    clear_w_x_4[2] = uSystolicPE_258_io_clear_w_d;
    clear_w_x_4[3] = uSystolicPE_273_io_clear_w_d;
    clear_w_x_4[4] = uSystolicPE_288_io_clear_w_d;
    clear_w_x_4[5] = uSystolicPE_303_io_clear_w_d;
    clear_w_x_4[6] = uSystolicPE_318_io_clear_w_d;
    clear_w_x_4[7] = uSystolicPE_333_io_clear_w_d;
    clear_w_x_4[8] = uSystolicPE_348_io_clear_w_d;
    clear_w_x_4[9] = uSystolicPE_363_io_clear_w_d;
    clear_w_x_4[10] = uSystolicPE_378_io_clear_w_d;
    clear_w_x_4[11] = uSystolicPE_393_io_clear_w_d;
    clear_w_x_4[12] = uSystolicPE_408_io_clear_w_d;
    clear_w_x_4[13] = uSystolicPE_423_io_clear_w_d;
    clear_w_x_4[14] = uSystolicPE_438_io_clear_w_d;
    clear_w_x_4[15] = uSystolicPE_453_io_clear_w_d;
    clear_w_x_4[16] = uSystolicPE_468_io_clear_w_d;
  end

  assign wght_sign_x_4_0 = io_wght_sign[4];
  assign wght_abs_x_4_0 = io_wght_abs_4;
  always @(*) begin
    enable_o_x_4[16] = io_enable_o[4];
    enable_o_x_4[0] = uSystolicPE_243_io_enable_o_d;
    enable_o_x_4[1] = uSystolicPE_258_io_enable_o_d;
    enable_o_x_4[2] = uSystolicPE_273_io_enable_o_d;
    enable_o_x_4[3] = uSystolicPE_288_io_enable_o_d;
    enable_o_x_4[4] = uSystolicPE_303_io_enable_o_d;
    enable_o_x_4[5] = uSystolicPE_318_io_enable_o_d;
    enable_o_x_4[6] = uSystolicPE_333_io_enable_o_d;
    enable_o_x_4[7] = uSystolicPE_348_io_enable_o_d;
    enable_o_x_4[8] = uSystolicPE_363_io_enable_o_d;
    enable_o_x_4[9] = uSystolicPE_378_io_enable_o_d;
    enable_o_x_4[10] = uSystolicPE_393_io_enable_o_d;
    enable_o_x_4[11] = uSystolicPE_408_io_enable_o_d;
    enable_o_x_4[12] = uSystolicPE_423_io_enable_o_d;
    enable_o_x_4[13] = uSystolicPE_438_io_enable_o_d;
    enable_o_x_4[14] = uSystolicPE_453_io_enable_o_d;
    enable_o_x_4[15] = uSystolicPE_468_io_enable_o_d;
  end

  always @(*) begin
    clear_o_x_4[16] = io_clear_o[4];
    clear_o_x_4[0] = uSystolicPE_243_io_clear_o_d;
    clear_o_x_4[1] = uSystolicPE_258_io_clear_o_d;
    clear_o_x_4[2] = uSystolicPE_273_io_clear_o_d;
    clear_o_x_4[3] = uSystolicPE_288_io_clear_o_d;
    clear_o_x_4[4] = uSystolicPE_303_io_clear_o_d;
    clear_o_x_4[5] = uSystolicPE_318_io_clear_o_d;
    clear_o_x_4[6] = uSystolicPE_333_io_clear_o_d;
    clear_o_x_4[7] = uSystolicPE_348_io_clear_o_d;
    clear_o_x_4[8] = uSystolicPE_363_io_clear_o_d;
    clear_o_x_4[9] = uSystolicPE_378_io_clear_o_d;
    clear_o_x_4[10] = uSystolicPE_393_io_clear_o_d;
    clear_o_x_4[11] = uSystolicPE_408_io_clear_o_d;
    clear_o_x_4[12] = uSystolicPE_423_io_clear_o_d;
    clear_o_x_4[13] = uSystolicPE_438_io_clear_o_d;
    clear_o_x_4[14] = uSystolicPE_453_io_clear_o_d;
    clear_o_x_4[15] = uSystolicPE_468_io_clear_o_d;
  end

  assign io_ofm_4 = ofm_x_4_0;
  assign ofm_x_4_16 = 32'h00000000;
  always @(*) begin
    enable_i_x_5[0] = io_enable_i[5];
    enable_i_x_5[1] = uSystolicPEBorder_21_io_enable_i_d;
    enable_i_x_5[2] = uSystolicPE_315_io_enable_i_d;
    enable_i_x_5[3] = uSystolicPE_316_io_enable_i_d;
    enable_i_x_5[4] = uSystolicPE_317_io_enable_i_d;
    enable_i_x_5[5] = uSystolicPE_318_io_enable_i_d;
    enable_i_x_5[6] = uSystolicPE_319_io_enable_i_d;
    enable_i_x_5[7] = uSystolicPE_320_io_enable_i_d;
    enable_i_x_5[8] = uSystolicPE_321_io_enable_i_d;
    enable_i_x_5[9] = uSystolicPE_322_io_enable_i_d;
    enable_i_x_5[10] = uSystolicPE_323_io_enable_i_d;
    enable_i_x_5[11] = uSystolicPE_324_io_enable_i_d;
    enable_i_x_5[12] = uSystolicPE_325_io_enable_i_d;
    enable_i_x_5[13] = uSystolicPE_326_io_enable_i_d;
    enable_i_x_5[14] = uSystolicPE_327_io_enable_i_d;
    enable_i_x_5[15] = uSystolicPE_328_io_enable_i_d;
    enable_i_x_5[16] = uSystolicPE_329_io_enable_i_d;
  end

  always @(*) begin
    clear_i_x_5[0] = io_clear_i[5];
    clear_i_x_5[1] = uSystolicPEBorder_21_io_clear_i_d;
    clear_i_x_5[2] = uSystolicPE_315_io_clear_i_d;
    clear_i_x_5[3] = uSystolicPE_316_io_clear_i_d;
    clear_i_x_5[4] = uSystolicPE_317_io_clear_i_d;
    clear_i_x_5[5] = uSystolicPE_318_io_clear_i_d;
    clear_i_x_5[6] = uSystolicPE_319_io_clear_i_d;
    clear_i_x_5[7] = uSystolicPE_320_io_clear_i_d;
    clear_i_x_5[8] = uSystolicPE_321_io_clear_i_d;
    clear_i_x_5[9] = uSystolicPE_322_io_clear_i_d;
    clear_i_x_5[10] = uSystolicPE_323_io_clear_i_d;
    clear_i_x_5[11] = uSystolicPE_324_io_clear_i_d;
    clear_i_x_5[12] = uSystolicPE_325_io_clear_i_d;
    clear_i_x_5[13] = uSystolicPE_326_io_clear_i_d;
    clear_i_x_5[14] = uSystolicPE_327_io_clear_i_d;
    clear_i_x_5[15] = uSystolicPE_328_io_clear_i_d;
    clear_i_x_5[16] = uSystolicPE_329_io_clear_i_d;
  end

  always @(*) begin
    mac_done_x_5[0] = io_mac_done[5];
    mac_done_x_5[1] = uSystolicPEBorder_21_io_mac_done_d;
    mac_done_x_5[2] = uSystolicPE_315_io_mac_done_d;
    mac_done_x_5[3] = uSystolicPE_316_io_mac_done_d;
    mac_done_x_5[4] = uSystolicPE_317_io_mac_done_d;
    mac_done_x_5[5] = uSystolicPE_318_io_mac_done_d;
    mac_done_x_5[6] = uSystolicPE_319_io_mac_done_d;
    mac_done_x_5[7] = uSystolicPE_320_io_mac_done_d;
    mac_done_x_5[8] = uSystolicPE_321_io_mac_done_d;
    mac_done_x_5[9] = uSystolicPE_322_io_mac_done_d;
    mac_done_x_5[10] = uSystolicPE_323_io_mac_done_d;
    mac_done_x_5[11] = uSystolicPE_324_io_mac_done_d;
    mac_done_x_5[12] = uSystolicPE_325_io_mac_done_d;
    mac_done_x_5[13] = uSystolicPE_326_io_mac_done_d;
    mac_done_x_5[14] = uSystolicPE_327_io_mac_done_d;
    mac_done_x_5[15] = uSystolicPE_328_io_mac_done_d;
    mac_done_x_5[16] = uSystolicPE_329_io_mac_done_d;
  end

  always @(*) begin
    enable_w_x_5[0] = io_enable_w[5];
    enable_w_x_5[1] = uSystolicPE_244_io_enable_w_d;
    enable_w_x_5[2] = uSystolicPE_259_io_enable_w_d;
    enable_w_x_5[3] = uSystolicPE_274_io_enable_w_d;
    enable_w_x_5[4] = uSystolicPE_289_io_enable_w_d;
    enable_w_x_5[5] = uSystolicPE_304_io_enable_w_d;
    enable_w_x_5[6] = uSystolicPE_319_io_enable_w_d;
    enable_w_x_5[7] = uSystolicPE_334_io_enable_w_d;
    enable_w_x_5[8] = uSystolicPE_349_io_enable_w_d;
    enable_w_x_5[9] = uSystolicPE_364_io_enable_w_d;
    enable_w_x_5[10] = uSystolicPE_379_io_enable_w_d;
    enable_w_x_5[11] = uSystolicPE_394_io_enable_w_d;
    enable_w_x_5[12] = uSystolicPE_409_io_enable_w_d;
    enable_w_x_5[13] = uSystolicPE_424_io_enable_w_d;
    enable_w_x_5[14] = uSystolicPE_439_io_enable_w_d;
    enable_w_x_5[15] = uSystolicPE_454_io_enable_w_d;
    enable_w_x_5[16] = uSystolicPE_469_io_enable_w_d;
  end

  always @(*) begin
    clear_w_x_5[0] = io_clear_w[5];
    clear_w_x_5[1] = uSystolicPE_244_io_clear_w_d;
    clear_w_x_5[2] = uSystolicPE_259_io_clear_w_d;
    clear_w_x_5[3] = uSystolicPE_274_io_clear_w_d;
    clear_w_x_5[4] = uSystolicPE_289_io_clear_w_d;
    clear_w_x_5[5] = uSystolicPE_304_io_clear_w_d;
    clear_w_x_5[6] = uSystolicPE_319_io_clear_w_d;
    clear_w_x_5[7] = uSystolicPE_334_io_clear_w_d;
    clear_w_x_5[8] = uSystolicPE_349_io_clear_w_d;
    clear_w_x_5[9] = uSystolicPE_364_io_clear_w_d;
    clear_w_x_5[10] = uSystolicPE_379_io_clear_w_d;
    clear_w_x_5[11] = uSystolicPE_394_io_clear_w_d;
    clear_w_x_5[12] = uSystolicPE_409_io_clear_w_d;
    clear_w_x_5[13] = uSystolicPE_424_io_clear_w_d;
    clear_w_x_5[14] = uSystolicPE_439_io_clear_w_d;
    clear_w_x_5[15] = uSystolicPE_454_io_clear_w_d;
    clear_w_x_5[16] = uSystolicPE_469_io_clear_w_d;
  end

  assign wght_sign_x_5_0 = io_wght_sign[5];
  assign wght_abs_x_5_0 = io_wght_abs_5;
  always @(*) begin
    enable_o_x_5[16] = io_enable_o[5];
    enable_o_x_5[0] = uSystolicPE_244_io_enable_o_d;
    enable_o_x_5[1] = uSystolicPE_259_io_enable_o_d;
    enable_o_x_5[2] = uSystolicPE_274_io_enable_o_d;
    enable_o_x_5[3] = uSystolicPE_289_io_enable_o_d;
    enable_o_x_5[4] = uSystolicPE_304_io_enable_o_d;
    enable_o_x_5[5] = uSystolicPE_319_io_enable_o_d;
    enable_o_x_5[6] = uSystolicPE_334_io_enable_o_d;
    enable_o_x_5[7] = uSystolicPE_349_io_enable_o_d;
    enable_o_x_5[8] = uSystolicPE_364_io_enable_o_d;
    enable_o_x_5[9] = uSystolicPE_379_io_enable_o_d;
    enable_o_x_5[10] = uSystolicPE_394_io_enable_o_d;
    enable_o_x_5[11] = uSystolicPE_409_io_enable_o_d;
    enable_o_x_5[12] = uSystolicPE_424_io_enable_o_d;
    enable_o_x_5[13] = uSystolicPE_439_io_enable_o_d;
    enable_o_x_5[14] = uSystolicPE_454_io_enable_o_d;
    enable_o_x_5[15] = uSystolicPE_469_io_enable_o_d;
  end

  always @(*) begin
    clear_o_x_5[16] = io_clear_o[5];
    clear_o_x_5[0] = uSystolicPE_244_io_clear_o_d;
    clear_o_x_5[1] = uSystolicPE_259_io_clear_o_d;
    clear_o_x_5[2] = uSystolicPE_274_io_clear_o_d;
    clear_o_x_5[3] = uSystolicPE_289_io_clear_o_d;
    clear_o_x_5[4] = uSystolicPE_304_io_clear_o_d;
    clear_o_x_5[5] = uSystolicPE_319_io_clear_o_d;
    clear_o_x_5[6] = uSystolicPE_334_io_clear_o_d;
    clear_o_x_5[7] = uSystolicPE_349_io_clear_o_d;
    clear_o_x_5[8] = uSystolicPE_364_io_clear_o_d;
    clear_o_x_5[9] = uSystolicPE_379_io_clear_o_d;
    clear_o_x_5[10] = uSystolicPE_394_io_clear_o_d;
    clear_o_x_5[11] = uSystolicPE_409_io_clear_o_d;
    clear_o_x_5[12] = uSystolicPE_424_io_clear_o_d;
    clear_o_x_5[13] = uSystolicPE_439_io_clear_o_d;
    clear_o_x_5[14] = uSystolicPE_454_io_clear_o_d;
    clear_o_x_5[15] = uSystolicPE_469_io_clear_o_d;
  end

  assign io_ofm_5 = ofm_x_5_0;
  assign ofm_x_5_16 = 32'h00000000;
  always @(*) begin
    enable_i_x_6[0] = io_enable_i[6];
    enable_i_x_6[1] = uSystolicPEBorder_22_io_enable_i_d;
    enable_i_x_6[2] = uSystolicPE_330_io_enable_i_d;
    enable_i_x_6[3] = uSystolicPE_331_io_enable_i_d;
    enable_i_x_6[4] = uSystolicPE_332_io_enable_i_d;
    enable_i_x_6[5] = uSystolicPE_333_io_enable_i_d;
    enable_i_x_6[6] = uSystolicPE_334_io_enable_i_d;
    enable_i_x_6[7] = uSystolicPE_335_io_enable_i_d;
    enable_i_x_6[8] = uSystolicPE_336_io_enable_i_d;
    enable_i_x_6[9] = uSystolicPE_337_io_enable_i_d;
    enable_i_x_6[10] = uSystolicPE_338_io_enable_i_d;
    enable_i_x_6[11] = uSystolicPE_339_io_enable_i_d;
    enable_i_x_6[12] = uSystolicPE_340_io_enable_i_d;
    enable_i_x_6[13] = uSystolicPE_341_io_enable_i_d;
    enable_i_x_6[14] = uSystolicPE_342_io_enable_i_d;
    enable_i_x_6[15] = uSystolicPE_343_io_enable_i_d;
    enable_i_x_6[16] = uSystolicPE_344_io_enable_i_d;
  end

  always @(*) begin
    clear_i_x_6[0] = io_clear_i[6];
    clear_i_x_6[1] = uSystolicPEBorder_22_io_clear_i_d;
    clear_i_x_6[2] = uSystolicPE_330_io_clear_i_d;
    clear_i_x_6[3] = uSystolicPE_331_io_clear_i_d;
    clear_i_x_6[4] = uSystolicPE_332_io_clear_i_d;
    clear_i_x_6[5] = uSystolicPE_333_io_clear_i_d;
    clear_i_x_6[6] = uSystolicPE_334_io_clear_i_d;
    clear_i_x_6[7] = uSystolicPE_335_io_clear_i_d;
    clear_i_x_6[8] = uSystolicPE_336_io_clear_i_d;
    clear_i_x_6[9] = uSystolicPE_337_io_clear_i_d;
    clear_i_x_6[10] = uSystolicPE_338_io_clear_i_d;
    clear_i_x_6[11] = uSystolicPE_339_io_clear_i_d;
    clear_i_x_6[12] = uSystolicPE_340_io_clear_i_d;
    clear_i_x_6[13] = uSystolicPE_341_io_clear_i_d;
    clear_i_x_6[14] = uSystolicPE_342_io_clear_i_d;
    clear_i_x_6[15] = uSystolicPE_343_io_clear_i_d;
    clear_i_x_6[16] = uSystolicPE_344_io_clear_i_d;
  end

  always @(*) begin
    mac_done_x_6[0] = io_mac_done[6];
    mac_done_x_6[1] = uSystolicPEBorder_22_io_mac_done_d;
    mac_done_x_6[2] = uSystolicPE_330_io_mac_done_d;
    mac_done_x_6[3] = uSystolicPE_331_io_mac_done_d;
    mac_done_x_6[4] = uSystolicPE_332_io_mac_done_d;
    mac_done_x_6[5] = uSystolicPE_333_io_mac_done_d;
    mac_done_x_6[6] = uSystolicPE_334_io_mac_done_d;
    mac_done_x_6[7] = uSystolicPE_335_io_mac_done_d;
    mac_done_x_6[8] = uSystolicPE_336_io_mac_done_d;
    mac_done_x_6[9] = uSystolicPE_337_io_mac_done_d;
    mac_done_x_6[10] = uSystolicPE_338_io_mac_done_d;
    mac_done_x_6[11] = uSystolicPE_339_io_mac_done_d;
    mac_done_x_6[12] = uSystolicPE_340_io_mac_done_d;
    mac_done_x_6[13] = uSystolicPE_341_io_mac_done_d;
    mac_done_x_6[14] = uSystolicPE_342_io_mac_done_d;
    mac_done_x_6[15] = uSystolicPE_343_io_mac_done_d;
    mac_done_x_6[16] = uSystolicPE_344_io_mac_done_d;
  end

  always @(*) begin
    enable_w_x_6[0] = io_enable_w[6];
    enable_w_x_6[1] = uSystolicPE_245_io_enable_w_d;
    enable_w_x_6[2] = uSystolicPE_260_io_enable_w_d;
    enable_w_x_6[3] = uSystolicPE_275_io_enable_w_d;
    enable_w_x_6[4] = uSystolicPE_290_io_enable_w_d;
    enable_w_x_6[5] = uSystolicPE_305_io_enable_w_d;
    enable_w_x_6[6] = uSystolicPE_320_io_enable_w_d;
    enable_w_x_6[7] = uSystolicPE_335_io_enable_w_d;
    enable_w_x_6[8] = uSystolicPE_350_io_enable_w_d;
    enable_w_x_6[9] = uSystolicPE_365_io_enable_w_d;
    enable_w_x_6[10] = uSystolicPE_380_io_enable_w_d;
    enable_w_x_6[11] = uSystolicPE_395_io_enable_w_d;
    enable_w_x_6[12] = uSystolicPE_410_io_enable_w_d;
    enable_w_x_6[13] = uSystolicPE_425_io_enable_w_d;
    enable_w_x_6[14] = uSystolicPE_440_io_enable_w_d;
    enable_w_x_6[15] = uSystolicPE_455_io_enable_w_d;
    enable_w_x_6[16] = uSystolicPE_470_io_enable_w_d;
  end

  always @(*) begin
    clear_w_x_6[0] = io_clear_w[6];
    clear_w_x_6[1] = uSystolicPE_245_io_clear_w_d;
    clear_w_x_6[2] = uSystolicPE_260_io_clear_w_d;
    clear_w_x_6[3] = uSystolicPE_275_io_clear_w_d;
    clear_w_x_6[4] = uSystolicPE_290_io_clear_w_d;
    clear_w_x_6[5] = uSystolicPE_305_io_clear_w_d;
    clear_w_x_6[6] = uSystolicPE_320_io_clear_w_d;
    clear_w_x_6[7] = uSystolicPE_335_io_clear_w_d;
    clear_w_x_6[8] = uSystolicPE_350_io_clear_w_d;
    clear_w_x_6[9] = uSystolicPE_365_io_clear_w_d;
    clear_w_x_6[10] = uSystolicPE_380_io_clear_w_d;
    clear_w_x_6[11] = uSystolicPE_395_io_clear_w_d;
    clear_w_x_6[12] = uSystolicPE_410_io_clear_w_d;
    clear_w_x_6[13] = uSystolicPE_425_io_clear_w_d;
    clear_w_x_6[14] = uSystolicPE_440_io_clear_w_d;
    clear_w_x_6[15] = uSystolicPE_455_io_clear_w_d;
    clear_w_x_6[16] = uSystolicPE_470_io_clear_w_d;
  end

  assign wght_sign_x_6_0 = io_wght_sign[6];
  assign wght_abs_x_6_0 = io_wght_abs_6;
  always @(*) begin
    enable_o_x_6[16] = io_enable_o[6];
    enable_o_x_6[0] = uSystolicPE_245_io_enable_o_d;
    enable_o_x_6[1] = uSystolicPE_260_io_enable_o_d;
    enable_o_x_6[2] = uSystolicPE_275_io_enable_o_d;
    enable_o_x_6[3] = uSystolicPE_290_io_enable_o_d;
    enable_o_x_6[4] = uSystolicPE_305_io_enable_o_d;
    enable_o_x_6[5] = uSystolicPE_320_io_enable_o_d;
    enable_o_x_6[6] = uSystolicPE_335_io_enable_o_d;
    enable_o_x_6[7] = uSystolicPE_350_io_enable_o_d;
    enable_o_x_6[8] = uSystolicPE_365_io_enable_o_d;
    enable_o_x_6[9] = uSystolicPE_380_io_enable_o_d;
    enable_o_x_6[10] = uSystolicPE_395_io_enable_o_d;
    enable_o_x_6[11] = uSystolicPE_410_io_enable_o_d;
    enable_o_x_6[12] = uSystolicPE_425_io_enable_o_d;
    enable_o_x_6[13] = uSystolicPE_440_io_enable_o_d;
    enable_o_x_6[14] = uSystolicPE_455_io_enable_o_d;
    enable_o_x_6[15] = uSystolicPE_470_io_enable_o_d;
  end

  always @(*) begin
    clear_o_x_6[16] = io_clear_o[6];
    clear_o_x_6[0] = uSystolicPE_245_io_clear_o_d;
    clear_o_x_6[1] = uSystolicPE_260_io_clear_o_d;
    clear_o_x_6[2] = uSystolicPE_275_io_clear_o_d;
    clear_o_x_6[3] = uSystolicPE_290_io_clear_o_d;
    clear_o_x_6[4] = uSystolicPE_305_io_clear_o_d;
    clear_o_x_6[5] = uSystolicPE_320_io_clear_o_d;
    clear_o_x_6[6] = uSystolicPE_335_io_clear_o_d;
    clear_o_x_6[7] = uSystolicPE_350_io_clear_o_d;
    clear_o_x_6[8] = uSystolicPE_365_io_clear_o_d;
    clear_o_x_6[9] = uSystolicPE_380_io_clear_o_d;
    clear_o_x_6[10] = uSystolicPE_395_io_clear_o_d;
    clear_o_x_6[11] = uSystolicPE_410_io_clear_o_d;
    clear_o_x_6[12] = uSystolicPE_425_io_clear_o_d;
    clear_o_x_6[13] = uSystolicPE_440_io_clear_o_d;
    clear_o_x_6[14] = uSystolicPE_455_io_clear_o_d;
    clear_o_x_6[15] = uSystolicPE_470_io_clear_o_d;
  end

  assign io_ofm_6 = ofm_x_6_0;
  assign ofm_x_6_16 = 32'h00000000;
  always @(*) begin
    enable_i_x_7[0] = io_enable_i[7];
    enable_i_x_7[1] = uSystolicPEBorder_23_io_enable_i_d;
    enable_i_x_7[2] = uSystolicPE_345_io_enable_i_d;
    enable_i_x_7[3] = uSystolicPE_346_io_enable_i_d;
    enable_i_x_7[4] = uSystolicPE_347_io_enable_i_d;
    enable_i_x_7[5] = uSystolicPE_348_io_enable_i_d;
    enable_i_x_7[6] = uSystolicPE_349_io_enable_i_d;
    enable_i_x_7[7] = uSystolicPE_350_io_enable_i_d;
    enable_i_x_7[8] = uSystolicPE_351_io_enable_i_d;
    enable_i_x_7[9] = uSystolicPE_352_io_enable_i_d;
    enable_i_x_7[10] = uSystolicPE_353_io_enable_i_d;
    enable_i_x_7[11] = uSystolicPE_354_io_enable_i_d;
    enable_i_x_7[12] = uSystolicPE_355_io_enable_i_d;
    enable_i_x_7[13] = uSystolicPE_356_io_enable_i_d;
    enable_i_x_7[14] = uSystolicPE_357_io_enable_i_d;
    enable_i_x_7[15] = uSystolicPE_358_io_enable_i_d;
    enable_i_x_7[16] = uSystolicPE_359_io_enable_i_d;
  end

  always @(*) begin
    clear_i_x_7[0] = io_clear_i[7];
    clear_i_x_7[1] = uSystolicPEBorder_23_io_clear_i_d;
    clear_i_x_7[2] = uSystolicPE_345_io_clear_i_d;
    clear_i_x_7[3] = uSystolicPE_346_io_clear_i_d;
    clear_i_x_7[4] = uSystolicPE_347_io_clear_i_d;
    clear_i_x_7[5] = uSystolicPE_348_io_clear_i_d;
    clear_i_x_7[6] = uSystolicPE_349_io_clear_i_d;
    clear_i_x_7[7] = uSystolicPE_350_io_clear_i_d;
    clear_i_x_7[8] = uSystolicPE_351_io_clear_i_d;
    clear_i_x_7[9] = uSystolicPE_352_io_clear_i_d;
    clear_i_x_7[10] = uSystolicPE_353_io_clear_i_d;
    clear_i_x_7[11] = uSystolicPE_354_io_clear_i_d;
    clear_i_x_7[12] = uSystolicPE_355_io_clear_i_d;
    clear_i_x_7[13] = uSystolicPE_356_io_clear_i_d;
    clear_i_x_7[14] = uSystolicPE_357_io_clear_i_d;
    clear_i_x_7[15] = uSystolicPE_358_io_clear_i_d;
    clear_i_x_7[16] = uSystolicPE_359_io_clear_i_d;
  end

  always @(*) begin
    mac_done_x_7[0] = io_mac_done[7];
    mac_done_x_7[1] = uSystolicPEBorder_23_io_mac_done_d;
    mac_done_x_7[2] = uSystolicPE_345_io_mac_done_d;
    mac_done_x_7[3] = uSystolicPE_346_io_mac_done_d;
    mac_done_x_7[4] = uSystolicPE_347_io_mac_done_d;
    mac_done_x_7[5] = uSystolicPE_348_io_mac_done_d;
    mac_done_x_7[6] = uSystolicPE_349_io_mac_done_d;
    mac_done_x_7[7] = uSystolicPE_350_io_mac_done_d;
    mac_done_x_7[8] = uSystolicPE_351_io_mac_done_d;
    mac_done_x_7[9] = uSystolicPE_352_io_mac_done_d;
    mac_done_x_7[10] = uSystolicPE_353_io_mac_done_d;
    mac_done_x_7[11] = uSystolicPE_354_io_mac_done_d;
    mac_done_x_7[12] = uSystolicPE_355_io_mac_done_d;
    mac_done_x_7[13] = uSystolicPE_356_io_mac_done_d;
    mac_done_x_7[14] = uSystolicPE_357_io_mac_done_d;
    mac_done_x_7[15] = uSystolicPE_358_io_mac_done_d;
    mac_done_x_7[16] = uSystolicPE_359_io_mac_done_d;
  end

  always @(*) begin
    enable_w_x_7[0] = io_enable_w[7];
    enable_w_x_7[1] = uSystolicPE_246_io_enable_w_d;
    enable_w_x_7[2] = uSystolicPE_261_io_enable_w_d;
    enable_w_x_7[3] = uSystolicPE_276_io_enable_w_d;
    enable_w_x_7[4] = uSystolicPE_291_io_enable_w_d;
    enable_w_x_7[5] = uSystolicPE_306_io_enable_w_d;
    enable_w_x_7[6] = uSystolicPE_321_io_enable_w_d;
    enable_w_x_7[7] = uSystolicPE_336_io_enable_w_d;
    enable_w_x_7[8] = uSystolicPE_351_io_enable_w_d;
    enable_w_x_7[9] = uSystolicPE_366_io_enable_w_d;
    enable_w_x_7[10] = uSystolicPE_381_io_enable_w_d;
    enable_w_x_7[11] = uSystolicPE_396_io_enable_w_d;
    enable_w_x_7[12] = uSystolicPE_411_io_enable_w_d;
    enable_w_x_7[13] = uSystolicPE_426_io_enable_w_d;
    enable_w_x_7[14] = uSystolicPE_441_io_enable_w_d;
    enable_w_x_7[15] = uSystolicPE_456_io_enable_w_d;
    enable_w_x_7[16] = uSystolicPE_471_io_enable_w_d;
  end

  always @(*) begin
    clear_w_x_7[0] = io_clear_w[7];
    clear_w_x_7[1] = uSystolicPE_246_io_clear_w_d;
    clear_w_x_7[2] = uSystolicPE_261_io_clear_w_d;
    clear_w_x_7[3] = uSystolicPE_276_io_clear_w_d;
    clear_w_x_7[4] = uSystolicPE_291_io_clear_w_d;
    clear_w_x_7[5] = uSystolicPE_306_io_clear_w_d;
    clear_w_x_7[6] = uSystolicPE_321_io_clear_w_d;
    clear_w_x_7[7] = uSystolicPE_336_io_clear_w_d;
    clear_w_x_7[8] = uSystolicPE_351_io_clear_w_d;
    clear_w_x_7[9] = uSystolicPE_366_io_clear_w_d;
    clear_w_x_7[10] = uSystolicPE_381_io_clear_w_d;
    clear_w_x_7[11] = uSystolicPE_396_io_clear_w_d;
    clear_w_x_7[12] = uSystolicPE_411_io_clear_w_d;
    clear_w_x_7[13] = uSystolicPE_426_io_clear_w_d;
    clear_w_x_7[14] = uSystolicPE_441_io_clear_w_d;
    clear_w_x_7[15] = uSystolicPE_456_io_clear_w_d;
    clear_w_x_7[16] = uSystolicPE_471_io_clear_w_d;
  end

  assign wght_sign_x_7_0 = io_wght_sign[7];
  assign wght_abs_x_7_0 = io_wght_abs_7;
  always @(*) begin
    enable_o_x_7[16] = io_enable_o[7];
    enable_o_x_7[0] = uSystolicPE_246_io_enable_o_d;
    enable_o_x_7[1] = uSystolicPE_261_io_enable_o_d;
    enable_o_x_7[2] = uSystolicPE_276_io_enable_o_d;
    enable_o_x_7[3] = uSystolicPE_291_io_enable_o_d;
    enable_o_x_7[4] = uSystolicPE_306_io_enable_o_d;
    enable_o_x_7[5] = uSystolicPE_321_io_enable_o_d;
    enable_o_x_7[6] = uSystolicPE_336_io_enable_o_d;
    enable_o_x_7[7] = uSystolicPE_351_io_enable_o_d;
    enable_o_x_7[8] = uSystolicPE_366_io_enable_o_d;
    enable_o_x_7[9] = uSystolicPE_381_io_enable_o_d;
    enable_o_x_7[10] = uSystolicPE_396_io_enable_o_d;
    enable_o_x_7[11] = uSystolicPE_411_io_enable_o_d;
    enable_o_x_7[12] = uSystolicPE_426_io_enable_o_d;
    enable_o_x_7[13] = uSystolicPE_441_io_enable_o_d;
    enable_o_x_7[14] = uSystolicPE_456_io_enable_o_d;
    enable_o_x_7[15] = uSystolicPE_471_io_enable_o_d;
  end

  always @(*) begin
    clear_o_x_7[16] = io_clear_o[7];
    clear_o_x_7[0] = uSystolicPE_246_io_clear_o_d;
    clear_o_x_7[1] = uSystolicPE_261_io_clear_o_d;
    clear_o_x_7[2] = uSystolicPE_276_io_clear_o_d;
    clear_o_x_7[3] = uSystolicPE_291_io_clear_o_d;
    clear_o_x_7[4] = uSystolicPE_306_io_clear_o_d;
    clear_o_x_7[5] = uSystolicPE_321_io_clear_o_d;
    clear_o_x_7[6] = uSystolicPE_336_io_clear_o_d;
    clear_o_x_7[7] = uSystolicPE_351_io_clear_o_d;
    clear_o_x_7[8] = uSystolicPE_366_io_clear_o_d;
    clear_o_x_7[9] = uSystolicPE_381_io_clear_o_d;
    clear_o_x_7[10] = uSystolicPE_396_io_clear_o_d;
    clear_o_x_7[11] = uSystolicPE_411_io_clear_o_d;
    clear_o_x_7[12] = uSystolicPE_426_io_clear_o_d;
    clear_o_x_7[13] = uSystolicPE_441_io_clear_o_d;
    clear_o_x_7[14] = uSystolicPE_456_io_clear_o_d;
    clear_o_x_7[15] = uSystolicPE_471_io_clear_o_d;
  end

  assign io_ofm_7 = ofm_x_7_0;
  assign ofm_x_7_16 = 32'h00000000;
  always @(*) begin
    enable_i_x_8[0] = io_enable_i[8];
    enable_i_x_8[1] = uSystolicPEBorder_24_io_enable_i_d;
    enable_i_x_8[2] = uSystolicPE_360_io_enable_i_d;
    enable_i_x_8[3] = uSystolicPE_361_io_enable_i_d;
    enable_i_x_8[4] = uSystolicPE_362_io_enable_i_d;
    enable_i_x_8[5] = uSystolicPE_363_io_enable_i_d;
    enable_i_x_8[6] = uSystolicPE_364_io_enable_i_d;
    enable_i_x_8[7] = uSystolicPE_365_io_enable_i_d;
    enable_i_x_8[8] = uSystolicPE_366_io_enable_i_d;
    enable_i_x_8[9] = uSystolicPE_367_io_enable_i_d;
    enable_i_x_8[10] = uSystolicPE_368_io_enable_i_d;
    enable_i_x_8[11] = uSystolicPE_369_io_enable_i_d;
    enable_i_x_8[12] = uSystolicPE_370_io_enable_i_d;
    enable_i_x_8[13] = uSystolicPE_371_io_enable_i_d;
    enable_i_x_8[14] = uSystolicPE_372_io_enable_i_d;
    enable_i_x_8[15] = uSystolicPE_373_io_enable_i_d;
    enable_i_x_8[16] = uSystolicPE_374_io_enable_i_d;
  end

  always @(*) begin
    clear_i_x_8[0] = io_clear_i[8];
    clear_i_x_8[1] = uSystolicPEBorder_24_io_clear_i_d;
    clear_i_x_8[2] = uSystolicPE_360_io_clear_i_d;
    clear_i_x_8[3] = uSystolicPE_361_io_clear_i_d;
    clear_i_x_8[4] = uSystolicPE_362_io_clear_i_d;
    clear_i_x_8[5] = uSystolicPE_363_io_clear_i_d;
    clear_i_x_8[6] = uSystolicPE_364_io_clear_i_d;
    clear_i_x_8[7] = uSystolicPE_365_io_clear_i_d;
    clear_i_x_8[8] = uSystolicPE_366_io_clear_i_d;
    clear_i_x_8[9] = uSystolicPE_367_io_clear_i_d;
    clear_i_x_8[10] = uSystolicPE_368_io_clear_i_d;
    clear_i_x_8[11] = uSystolicPE_369_io_clear_i_d;
    clear_i_x_8[12] = uSystolicPE_370_io_clear_i_d;
    clear_i_x_8[13] = uSystolicPE_371_io_clear_i_d;
    clear_i_x_8[14] = uSystolicPE_372_io_clear_i_d;
    clear_i_x_8[15] = uSystolicPE_373_io_clear_i_d;
    clear_i_x_8[16] = uSystolicPE_374_io_clear_i_d;
  end

  always @(*) begin
    mac_done_x_8[0] = io_mac_done[8];
    mac_done_x_8[1] = uSystolicPEBorder_24_io_mac_done_d;
    mac_done_x_8[2] = uSystolicPE_360_io_mac_done_d;
    mac_done_x_8[3] = uSystolicPE_361_io_mac_done_d;
    mac_done_x_8[4] = uSystolicPE_362_io_mac_done_d;
    mac_done_x_8[5] = uSystolicPE_363_io_mac_done_d;
    mac_done_x_8[6] = uSystolicPE_364_io_mac_done_d;
    mac_done_x_8[7] = uSystolicPE_365_io_mac_done_d;
    mac_done_x_8[8] = uSystolicPE_366_io_mac_done_d;
    mac_done_x_8[9] = uSystolicPE_367_io_mac_done_d;
    mac_done_x_8[10] = uSystolicPE_368_io_mac_done_d;
    mac_done_x_8[11] = uSystolicPE_369_io_mac_done_d;
    mac_done_x_8[12] = uSystolicPE_370_io_mac_done_d;
    mac_done_x_8[13] = uSystolicPE_371_io_mac_done_d;
    mac_done_x_8[14] = uSystolicPE_372_io_mac_done_d;
    mac_done_x_8[15] = uSystolicPE_373_io_mac_done_d;
    mac_done_x_8[16] = uSystolicPE_374_io_mac_done_d;
  end

  always @(*) begin
    enable_w_x_8[0] = io_enable_w[8];
    enable_w_x_8[1] = uSystolicPE_247_io_enable_w_d;
    enable_w_x_8[2] = uSystolicPE_262_io_enable_w_d;
    enable_w_x_8[3] = uSystolicPE_277_io_enable_w_d;
    enable_w_x_8[4] = uSystolicPE_292_io_enable_w_d;
    enable_w_x_8[5] = uSystolicPE_307_io_enable_w_d;
    enable_w_x_8[6] = uSystolicPE_322_io_enable_w_d;
    enable_w_x_8[7] = uSystolicPE_337_io_enable_w_d;
    enable_w_x_8[8] = uSystolicPE_352_io_enable_w_d;
    enable_w_x_8[9] = uSystolicPE_367_io_enable_w_d;
    enable_w_x_8[10] = uSystolicPE_382_io_enable_w_d;
    enable_w_x_8[11] = uSystolicPE_397_io_enable_w_d;
    enable_w_x_8[12] = uSystolicPE_412_io_enable_w_d;
    enable_w_x_8[13] = uSystolicPE_427_io_enable_w_d;
    enable_w_x_8[14] = uSystolicPE_442_io_enable_w_d;
    enable_w_x_8[15] = uSystolicPE_457_io_enable_w_d;
    enable_w_x_8[16] = uSystolicPE_472_io_enable_w_d;
  end

  always @(*) begin
    clear_w_x_8[0] = io_clear_w[8];
    clear_w_x_8[1] = uSystolicPE_247_io_clear_w_d;
    clear_w_x_8[2] = uSystolicPE_262_io_clear_w_d;
    clear_w_x_8[3] = uSystolicPE_277_io_clear_w_d;
    clear_w_x_8[4] = uSystolicPE_292_io_clear_w_d;
    clear_w_x_8[5] = uSystolicPE_307_io_clear_w_d;
    clear_w_x_8[6] = uSystolicPE_322_io_clear_w_d;
    clear_w_x_8[7] = uSystolicPE_337_io_clear_w_d;
    clear_w_x_8[8] = uSystolicPE_352_io_clear_w_d;
    clear_w_x_8[9] = uSystolicPE_367_io_clear_w_d;
    clear_w_x_8[10] = uSystolicPE_382_io_clear_w_d;
    clear_w_x_8[11] = uSystolicPE_397_io_clear_w_d;
    clear_w_x_8[12] = uSystolicPE_412_io_clear_w_d;
    clear_w_x_8[13] = uSystolicPE_427_io_clear_w_d;
    clear_w_x_8[14] = uSystolicPE_442_io_clear_w_d;
    clear_w_x_8[15] = uSystolicPE_457_io_clear_w_d;
    clear_w_x_8[16] = uSystolicPE_472_io_clear_w_d;
  end

  assign wght_sign_x_8_0 = io_wght_sign[8];
  assign wght_abs_x_8_0 = io_wght_abs_8;
  always @(*) begin
    enable_o_x_8[16] = io_enable_o[8];
    enable_o_x_8[0] = uSystolicPE_247_io_enable_o_d;
    enable_o_x_8[1] = uSystolicPE_262_io_enable_o_d;
    enable_o_x_8[2] = uSystolicPE_277_io_enable_o_d;
    enable_o_x_8[3] = uSystolicPE_292_io_enable_o_d;
    enable_o_x_8[4] = uSystolicPE_307_io_enable_o_d;
    enable_o_x_8[5] = uSystolicPE_322_io_enable_o_d;
    enable_o_x_8[6] = uSystolicPE_337_io_enable_o_d;
    enable_o_x_8[7] = uSystolicPE_352_io_enable_o_d;
    enable_o_x_8[8] = uSystolicPE_367_io_enable_o_d;
    enable_o_x_8[9] = uSystolicPE_382_io_enable_o_d;
    enable_o_x_8[10] = uSystolicPE_397_io_enable_o_d;
    enable_o_x_8[11] = uSystolicPE_412_io_enable_o_d;
    enable_o_x_8[12] = uSystolicPE_427_io_enable_o_d;
    enable_o_x_8[13] = uSystolicPE_442_io_enable_o_d;
    enable_o_x_8[14] = uSystolicPE_457_io_enable_o_d;
    enable_o_x_8[15] = uSystolicPE_472_io_enable_o_d;
  end

  always @(*) begin
    clear_o_x_8[16] = io_clear_o[8];
    clear_o_x_8[0] = uSystolicPE_247_io_clear_o_d;
    clear_o_x_8[1] = uSystolicPE_262_io_clear_o_d;
    clear_o_x_8[2] = uSystolicPE_277_io_clear_o_d;
    clear_o_x_8[3] = uSystolicPE_292_io_clear_o_d;
    clear_o_x_8[4] = uSystolicPE_307_io_clear_o_d;
    clear_o_x_8[5] = uSystolicPE_322_io_clear_o_d;
    clear_o_x_8[6] = uSystolicPE_337_io_clear_o_d;
    clear_o_x_8[7] = uSystolicPE_352_io_clear_o_d;
    clear_o_x_8[8] = uSystolicPE_367_io_clear_o_d;
    clear_o_x_8[9] = uSystolicPE_382_io_clear_o_d;
    clear_o_x_8[10] = uSystolicPE_397_io_clear_o_d;
    clear_o_x_8[11] = uSystolicPE_412_io_clear_o_d;
    clear_o_x_8[12] = uSystolicPE_427_io_clear_o_d;
    clear_o_x_8[13] = uSystolicPE_442_io_clear_o_d;
    clear_o_x_8[14] = uSystolicPE_457_io_clear_o_d;
    clear_o_x_8[15] = uSystolicPE_472_io_clear_o_d;
  end

  assign io_ofm_8 = ofm_x_8_0;
  assign ofm_x_8_16 = 32'h00000000;
  always @(*) begin
    enable_i_x_9[0] = io_enable_i[9];
    enable_i_x_9[1] = uSystolicPEBorder_25_io_enable_i_d;
    enable_i_x_9[2] = uSystolicPE_375_io_enable_i_d;
    enable_i_x_9[3] = uSystolicPE_376_io_enable_i_d;
    enable_i_x_9[4] = uSystolicPE_377_io_enable_i_d;
    enable_i_x_9[5] = uSystolicPE_378_io_enable_i_d;
    enable_i_x_9[6] = uSystolicPE_379_io_enable_i_d;
    enable_i_x_9[7] = uSystolicPE_380_io_enable_i_d;
    enable_i_x_9[8] = uSystolicPE_381_io_enable_i_d;
    enable_i_x_9[9] = uSystolicPE_382_io_enable_i_d;
    enable_i_x_9[10] = uSystolicPE_383_io_enable_i_d;
    enable_i_x_9[11] = uSystolicPE_384_io_enable_i_d;
    enable_i_x_9[12] = uSystolicPE_385_io_enable_i_d;
    enable_i_x_9[13] = uSystolicPE_386_io_enable_i_d;
    enable_i_x_9[14] = uSystolicPE_387_io_enable_i_d;
    enable_i_x_9[15] = uSystolicPE_388_io_enable_i_d;
    enable_i_x_9[16] = uSystolicPE_389_io_enable_i_d;
  end

  always @(*) begin
    clear_i_x_9[0] = io_clear_i[9];
    clear_i_x_9[1] = uSystolicPEBorder_25_io_clear_i_d;
    clear_i_x_9[2] = uSystolicPE_375_io_clear_i_d;
    clear_i_x_9[3] = uSystolicPE_376_io_clear_i_d;
    clear_i_x_9[4] = uSystolicPE_377_io_clear_i_d;
    clear_i_x_9[5] = uSystolicPE_378_io_clear_i_d;
    clear_i_x_9[6] = uSystolicPE_379_io_clear_i_d;
    clear_i_x_9[7] = uSystolicPE_380_io_clear_i_d;
    clear_i_x_9[8] = uSystolicPE_381_io_clear_i_d;
    clear_i_x_9[9] = uSystolicPE_382_io_clear_i_d;
    clear_i_x_9[10] = uSystolicPE_383_io_clear_i_d;
    clear_i_x_9[11] = uSystolicPE_384_io_clear_i_d;
    clear_i_x_9[12] = uSystolicPE_385_io_clear_i_d;
    clear_i_x_9[13] = uSystolicPE_386_io_clear_i_d;
    clear_i_x_9[14] = uSystolicPE_387_io_clear_i_d;
    clear_i_x_9[15] = uSystolicPE_388_io_clear_i_d;
    clear_i_x_9[16] = uSystolicPE_389_io_clear_i_d;
  end

  always @(*) begin
    mac_done_x_9[0] = io_mac_done[9];
    mac_done_x_9[1] = uSystolicPEBorder_25_io_mac_done_d;
    mac_done_x_9[2] = uSystolicPE_375_io_mac_done_d;
    mac_done_x_9[3] = uSystolicPE_376_io_mac_done_d;
    mac_done_x_9[4] = uSystolicPE_377_io_mac_done_d;
    mac_done_x_9[5] = uSystolicPE_378_io_mac_done_d;
    mac_done_x_9[6] = uSystolicPE_379_io_mac_done_d;
    mac_done_x_9[7] = uSystolicPE_380_io_mac_done_d;
    mac_done_x_9[8] = uSystolicPE_381_io_mac_done_d;
    mac_done_x_9[9] = uSystolicPE_382_io_mac_done_d;
    mac_done_x_9[10] = uSystolicPE_383_io_mac_done_d;
    mac_done_x_9[11] = uSystolicPE_384_io_mac_done_d;
    mac_done_x_9[12] = uSystolicPE_385_io_mac_done_d;
    mac_done_x_9[13] = uSystolicPE_386_io_mac_done_d;
    mac_done_x_9[14] = uSystolicPE_387_io_mac_done_d;
    mac_done_x_9[15] = uSystolicPE_388_io_mac_done_d;
    mac_done_x_9[16] = uSystolicPE_389_io_mac_done_d;
  end

  always @(*) begin
    enable_w_x_9[0] = io_enable_w[9];
    enable_w_x_9[1] = uSystolicPE_248_io_enable_w_d;
    enable_w_x_9[2] = uSystolicPE_263_io_enable_w_d;
    enable_w_x_9[3] = uSystolicPE_278_io_enable_w_d;
    enable_w_x_9[4] = uSystolicPE_293_io_enable_w_d;
    enable_w_x_9[5] = uSystolicPE_308_io_enable_w_d;
    enable_w_x_9[6] = uSystolicPE_323_io_enable_w_d;
    enable_w_x_9[7] = uSystolicPE_338_io_enable_w_d;
    enable_w_x_9[8] = uSystolicPE_353_io_enable_w_d;
    enable_w_x_9[9] = uSystolicPE_368_io_enable_w_d;
    enable_w_x_9[10] = uSystolicPE_383_io_enable_w_d;
    enable_w_x_9[11] = uSystolicPE_398_io_enable_w_d;
    enable_w_x_9[12] = uSystolicPE_413_io_enable_w_d;
    enable_w_x_9[13] = uSystolicPE_428_io_enable_w_d;
    enable_w_x_9[14] = uSystolicPE_443_io_enable_w_d;
    enable_w_x_9[15] = uSystolicPE_458_io_enable_w_d;
    enable_w_x_9[16] = uSystolicPE_473_io_enable_w_d;
  end

  always @(*) begin
    clear_w_x_9[0] = io_clear_w[9];
    clear_w_x_9[1] = uSystolicPE_248_io_clear_w_d;
    clear_w_x_9[2] = uSystolicPE_263_io_clear_w_d;
    clear_w_x_9[3] = uSystolicPE_278_io_clear_w_d;
    clear_w_x_9[4] = uSystolicPE_293_io_clear_w_d;
    clear_w_x_9[5] = uSystolicPE_308_io_clear_w_d;
    clear_w_x_9[6] = uSystolicPE_323_io_clear_w_d;
    clear_w_x_9[7] = uSystolicPE_338_io_clear_w_d;
    clear_w_x_9[8] = uSystolicPE_353_io_clear_w_d;
    clear_w_x_9[9] = uSystolicPE_368_io_clear_w_d;
    clear_w_x_9[10] = uSystolicPE_383_io_clear_w_d;
    clear_w_x_9[11] = uSystolicPE_398_io_clear_w_d;
    clear_w_x_9[12] = uSystolicPE_413_io_clear_w_d;
    clear_w_x_9[13] = uSystolicPE_428_io_clear_w_d;
    clear_w_x_9[14] = uSystolicPE_443_io_clear_w_d;
    clear_w_x_9[15] = uSystolicPE_458_io_clear_w_d;
    clear_w_x_9[16] = uSystolicPE_473_io_clear_w_d;
  end

  assign wght_sign_x_9_0 = io_wght_sign[9];
  assign wght_abs_x_9_0 = io_wght_abs_9;
  always @(*) begin
    enable_o_x_9[16] = io_enable_o[9];
    enable_o_x_9[0] = uSystolicPE_248_io_enable_o_d;
    enable_o_x_9[1] = uSystolicPE_263_io_enable_o_d;
    enable_o_x_9[2] = uSystolicPE_278_io_enable_o_d;
    enable_o_x_9[3] = uSystolicPE_293_io_enable_o_d;
    enable_o_x_9[4] = uSystolicPE_308_io_enable_o_d;
    enable_o_x_9[5] = uSystolicPE_323_io_enable_o_d;
    enable_o_x_9[6] = uSystolicPE_338_io_enable_o_d;
    enable_o_x_9[7] = uSystolicPE_353_io_enable_o_d;
    enable_o_x_9[8] = uSystolicPE_368_io_enable_o_d;
    enable_o_x_9[9] = uSystolicPE_383_io_enable_o_d;
    enable_o_x_9[10] = uSystolicPE_398_io_enable_o_d;
    enable_o_x_9[11] = uSystolicPE_413_io_enable_o_d;
    enable_o_x_9[12] = uSystolicPE_428_io_enable_o_d;
    enable_o_x_9[13] = uSystolicPE_443_io_enable_o_d;
    enable_o_x_9[14] = uSystolicPE_458_io_enable_o_d;
    enable_o_x_9[15] = uSystolicPE_473_io_enable_o_d;
  end

  always @(*) begin
    clear_o_x_9[16] = io_clear_o[9];
    clear_o_x_9[0] = uSystolicPE_248_io_clear_o_d;
    clear_o_x_9[1] = uSystolicPE_263_io_clear_o_d;
    clear_o_x_9[2] = uSystolicPE_278_io_clear_o_d;
    clear_o_x_9[3] = uSystolicPE_293_io_clear_o_d;
    clear_o_x_9[4] = uSystolicPE_308_io_clear_o_d;
    clear_o_x_9[5] = uSystolicPE_323_io_clear_o_d;
    clear_o_x_9[6] = uSystolicPE_338_io_clear_o_d;
    clear_o_x_9[7] = uSystolicPE_353_io_clear_o_d;
    clear_o_x_9[8] = uSystolicPE_368_io_clear_o_d;
    clear_o_x_9[9] = uSystolicPE_383_io_clear_o_d;
    clear_o_x_9[10] = uSystolicPE_398_io_clear_o_d;
    clear_o_x_9[11] = uSystolicPE_413_io_clear_o_d;
    clear_o_x_9[12] = uSystolicPE_428_io_clear_o_d;
    clear_o_x_9[13] = uSystolicPE_443_io_clear_o_d;
    clear_o_x_9[14] = uSystolicPE_458_io_clear_o_d;
    clear_o_x_9[15] = uSystolicPE_473_io_clear_o_d;
  end

  assign io_ofm_9 = ofm_x_9_0;
  assign ofm_x_9_16 = 32'h00000000;
  always @(*) begin
    enable_i_x_10[0] = io_enable_i[10];
    enable_i_x_10[1] = uSystolicPEBorder_26_io_enable_i_d;
    enable_i_x_10[2] = uSystolicPE_390_io_enable_i_d;
    enable_i_x_10[3] = uSystolicPE_391_io_enable_i_d;
    enable_i_x_10[4] = uSystolicPE_392_io_enable_i_d;
    enable_i_x_10[5] = uSystolicPE_393_io_enable_i_d;
    enable_i_x_10[6] = uSystolicPE_394_io_enable_i_d;
    enable_i_x_10[7] = uSystolicPE_395_io_enable_i_d;
    enable_i_x_10[8] = uSystolicPE_396_io_enable_i_d;
    enable_i_x_10[9] = uSystolicPE_397_io_enable_i_d;
    enable_i_x_10[10] = uSystolicPE_398_io_enable_i_d;
    enable_i_x_10[11] = uSystolicPE_399_io_enable_i_d;
    enable_i_x_10[12] = uSystolicPE_400_io_enable_i_d;
    enable_i_x_10[13] = uSystolicPE_401_io_enable_i_d;
    enable_i_x_10[14] = uSystolicPE_402_io_enable_i_d;
    enable_i_x_10[15] = uSystolicPE_403_io_enable_i_d;
    enable_i_x_10[16] = uSystolicPE_404_io_enable_i_d;
  end

  always @(*) begin
    clear_i_x_10[0] = io_clear_i[10];
    clear_i_x_10[1] = uSystolicPEBorder_26_io_clear_i_d;
    clear_i_x_10[2] = uSystolicPE_390_io_clear_i_d;
    clear_i_x_10[3] = uSystolicPE_391_io_clear_i_d;
    clear_i_x_10[4] = uSystolicPE_392_io_clear_i_d;
    clear_i_x_10[5] = uSystolicPE_393_io_clear_i_d;
    clear_i_x_10[6] = uSystolicPE_394_io_clear_i_d;
    clear_i_x_10[7] = uSystolicPE_395_io_clear_i_d;
    clear_i_x_10[8] = uSystolicPE_396_io_clear_i_d;
    clear_i_x_10[9] = uSystolicPE_397_io_clear_i_d;
    clear_i_x_10[10] = uSystolicPE_398_io_clear_i_d;
    clear_i_x_10[11] = uSystolicPE_399_io_clear_i_d;
    clear_i_x_10[12] = uSystolicPE_400_io_clear_i_d;
    clear_i_x_10[13] = uSystolicPE_401_io_clear_i_d;
    clear_i_x_10[14] = uSystolicPE_402_io_clear_i_d;
    clear_i_x_10[15] = uSystolicPE_403_io_clear_i_d;
    clear_i_x_10[16] = uSystolicPE_404_io_clear_i_d;
  end

  always @(*) begin
    mac_done_x_10[0] = io_mac_done[10];
    mac_done_x_10[1] = uSystolicPEBorder_26_io_mac_done_d;
    mac_done_x_10[2] = uSystolicPE_390_io_mac_done_d;
    mac_done_x_10[3] = uSystolicPE_391_io_mac_done_d;
    mac_done_x_10[4] = uSystolicPE_392_io_mac_done_d;
    mac_done_x_10[5] = uSystolicPE_393_io_mac_done_d;
    mac_done_x_10[6] = uSystolicPE_394_io_mac_done_d;
    mac_done_x_10[7] = uSystolicPE_395_io_mac_done_d;
    mac_done_x_10[8] = uSystolicPE_396_io_mac_done_d;
    mac_done_x_10[9] = uSystolicPE_397_io_mac_done_d;
    mac_done_x_10[10] = uSystolicPE_398_io_mac_done_d;
    mac_done_x_10[11] = uSystolicPE_399_io_mac_done_d;
    mac_done_x_10[12] = uSystolicPE_400_io_mac_done_d;
    mac_done_x_10[13] = uSystolicPE_401_io_mac_done_d;
    mac_done_x_10[14] = uSystolicPE_402_io_mac_done_d;
    mac_done_x_10[15] = uSystolicPE_403_io_mac_done_d;
    mac_done_x_10[16] = uSystolicPE_404_io_mac_done_d;
  end

  always @(*) begin
    enable_w_x_10[0] = io_enable_w[10];
    enable_w_x_10[1] = uSystolicPE_249_io_enable_w_d;
    enable_w_x_10[2] = uSystolicPE_264_io_enable_w_d;
    enable_w_x_10[3] = uSystolicPE_279_io_enable_w_d;
    enable_w_x_10[4] = uSystolicPE_294_io_enable_w_d;
    enable_w_x_10[5] = uSystolicPE_309_io_enable_w_d;
    enable_w_x_10[6] = uSystolicPE_324_io_enable_w_d;
    enable_w_x_10[7] = uSystolicPE_339_io_enable_w_d;
    enable_w_x_10[8] = uSystolicPE_354_io_enable_w_d;
    enable_w_x_10[9] = uSystolicPE_369_io_enable_w_d;
    enable_w_x_10[10] = uSystolicPE_384_io_enable_w_d;
    enable_w_x_10[11] = uSystolicPE_399_io_enable_w_d;
    enable_w_x_10[12] = uSystolicPE_414_io_enable_w_d;
    enable_w_x_10[13] = uSystolicPE_429_io_enable_w_d;
    enable_w_x_10[14] = uSystolicPE_444_io_enable_w_d;
    enable_w_x_10[15] = uSystolicPE_459_io_enable_w_d;
    enable_w_x_10[16] = uSystolicPE_474_io_enable_w_d;
  end

  always @(*) begin
    clear_w_x_10[0] = io_clear_w[10];
    clear_w_x_10[1] = uSystolicPE_249_io_clear_w_d;
    clear_w_x_10[2] = uSystolicPE_264_io_clear_w_d;
    clear_w_x_10[3] = uSystolicPE_279_io_clear_w_d;
    clear_w_x_10[4] = uSystolicPE_294_io_clear_w_d;
    clear_w_x_10[5] = uSystolicPE_309_io_clear_w_d;
    clear_w_x_10[6] = uSystolicPE_324_io_clear_w_d;
    clear_w_x_10[7] = uSystolicPE_339_io_clear_w_d;
    clear_w_x_10[8] = uSystolicPE_354_io_clear_w_d;
    clear_w_x_10[9] = uSystolicPE_369_io_clear_w_d;
    clear_w_x_10[10] = uSystolicPE_384_io_clear_w_d;
    clear_w_x_10[11] = uSystolicPE_399_io_clear_w_d;
    clear_w_x_10[12] = uSystolicPE_414_io_clear_w_d;
    clear_w_x_10[13] = uSystolicPE_429_io_clear_w_d;
    clear_w_x_10[14] = uSystolicPE_444_io_clear_w_d;
    clear_w_x_10[15] = uSystolicPE_459_io_clear_w_d;
    clear_w_x_10[16] = uSystolicPE_474_io_clear_w_d;
  end

  assign wght_sign_x_10_0 = io_wght_sign[10];
  assign wght_abs_x_10_0 = io_wght_abs_10;
  always @(*) begin
    enable_o_x_10[16] = io_enable_o[10];
    enable_o_x_10[0] = uSystolicPE_249_io_enable_o_d;
    enable_o_x_10[1] = uSystolicPE_264_io_enable_o_d;
    enable_o_x_10[2] = uSystolicPE_279_io_enable_o_d;
    enable_o_x_10[3] = uSystolicPE_294_io_enable_o_d;
    enable_o_x_10[4] = uSystolicPE_309_io_enable_o_d;
    enable_o_x_10[5] = uSystolicPE_324_io_enable_o_d;
    enable_o_x_10[6] = uSystolicPE_339_io_enable_o_d;
    enable_o_x_10[7] = uSystolicPE_354_io_enable_o_d;
    enable_o_x_10[8] = uSystolicPE_369_io_enable_o_d;
    enable_o_x_10[9] = uSystolicPE_384_io_enable_o_d;
    enable_o_x_10[10] = uSystolicPE_399_io_enable_o_d;
    enable_o_x_10[11] = uSystolicPE_414_io_enable_o_d;
    enable_o_x_10[12] = uSystolicPE_429_io_enable_o_d;
    enable_o_x_10[13] = uSystolicPE_444_io_enable_o_d;
    enable_o_x_10[14] = uSystolicPE_459_io_enable_o_d;
    enable_o_x_10[15] = uSystolicPE_474_io_enable_o_d;
  end

  always @(*) begin
    clear_o_x_10[16] = io_clear_o[10];
    clear_o_x_10[0] = uSystolicPE_249_io_clear_o_d;
    clear_o_x_10[1] = uSystolicPE_264_io_clear_o_d;
    clear_o_x_10[2] = uSystolicPE_279_io_clear_o_d;
    clear_o_x_10[3] = uSystolicPE_294_io_clear_o_d;
    clear_o_x_10[4] = uSystolicPE_309_io_clear_o_d;
    clear_o_x_10[5] = uSystolicPE_324_io_clear_o_d;
    clear_o_x_10[6] = uSystolicPE_339_io_clear_o_d;
    clear_o_x_10[7] = uSystolicPE_354_io_clear_o_d;
    clear_o_x_10[8] = uSystolicPE_369_io_clear_o_d;
    clear_o_x_10[9] = uSystolicPE_384_io_clear_o_d;
    clear_o_x_10[10] = uSystolicPE_399_io_clear_o_d;
    clear_o_x_10[11] = uSystolicPE_414_io_clear_o_d;
    clear_o_x_10[12] = uSystolicPE_429_io_clear_o_d;
    clear_o_x_10[13] = uSystolicPE_444_io_clear_o_d;
    clear_o_x_10[14] = uSystolicPE_459_io_clear_o_d;
    clear_o_x_10[15] = uSystolicPE_474_io_clear_o_d;
  end

  assign io_ofm_10 = ofm_x_10_0;
  assign ofm_x_10_16 = 32'h00000000;
  always @(*) begin
    enable_i_x_11[0] = io_enable_i[11];
    enable_i_x_11[1] = uSystolicPEBorder_27_io_enable_i_d;
    enable_i_x_11[2] = uSystolicPE_405_io_enable_i_d;
    enable_i_x_11[3] = uSystolicPE_406_io_enable_i_d;
    enable_i_x_11[4] = uSystolicPE_407_io_enable_i_d;
    enable_i_x_11[5] = uSystolicPE_408_io_enable_i_d;
    enable_i_x_11[6] = uSystolicPE_409_io_enable_i_d;
    enable_i_x_11[7] = uSystolicPE_410_io_enable_i_d;
    enable_i_x_11[8] = uSystolicPE_411_io_enable_i_d;
    enable_i_x_11[9] = uSystolicPE_412_io_enable_i_d;
    enable_i_x_11[10] = uSystolicPE_413_io_enable_i_d;
    enable_i_x_11[11] = uSystolicPE_414_io_enable_i_d;
    enable_i_x_11[12] = uSystolicPE_415_io_enable_i_d;
    enable_i_x_11[13] = uSystolicPE_416_io_enable_i_d;
    enable_i_x_11[14] = uSystolicPE_417_io_enable_i_d;
    enable_i_x_11[15] = uSystolicPE_418_io_enable_i_d;
    enable_i_x_11[16] = uSystolicPE_419_io_enable_i_d;
  end

  always @(*) begin
    clear_i_x_11[0] = io_clear_i[11];
    clear_i_x_11[1] = uSystolicPEBorder_27_io_clear_i_d;
    clear_i_x_11[2] = uSystolicPE_405_io_clear_i_d;
    clear_i_x_11[3] = uSystolicPE_406_io_clear_i_d;
    clear_i_x_11[4] = uSystolicPE_407_io_clear_i_d;
    clear_i_x_11[5] = uSystolicPE_408_io_clear_i_d;
    clear_i_x_11[6] = uSystolicPE_409_io_clear_i_d;
    clear_i_x_11[7] = uSystolicPE_410_io_clear_i_d;
    clear_i_x_11[8] = uSystolicPE_411_io_clear_i_d;
    clear_i_x_11[9] = uSystolicPE_412_io_clear_i_d;
    clear_i_x_11[10] = uSystolicPE_413_io_clear_i_d;
    clear_i_x_11[11] = uSystolicPE_414_io_clear_i_d;
    clear_i_x_11[12] = uSystolicPE_415_io_clear_i_d;
    clear_i_x_11[13] = uSystolicPE_416_io_clear_i_d;
    clear_i_x_11[14] = uSystolicPE_417_io_clear_i_d;
    clear_i_x_11[15] = uSystolicPE_418_io_clear_i_d;
    clear_i_x_11[16] = uSystolicPE_419_io_clear_i_d;
  end

  always @(*) begin
    mac_done_x_11[0] = io_mac_done[11];
    mac_done_x_11[1] = uSystolicPEBorder_27_io_mac_done_d;
    mac_done_x_11[2] = uSystolicPE_405_io_mac_done_d;
    mac_done_x_11[3] = uSystolicPE_406_io_mac_done_d;
    mac_done_x_11[4] = uSystolicPE_407_io_mac_done_d;
    mac_done_x_11[5] = uSystolicPE_408_io_mac_done_d;
    mac_done_x_11[6] = uSystolicPE_409_io_mac_done_d;
    mac_done_x_11[7] = uSystolicPE_410_io_mac_done_d;
    mac_done_x_11[8] = uSystolicPE_411_io_mac_done_d;
    mac_done_x_11[9] = uSystolicPE_412_io_mac_done_d;
    mac_done_x_11[10] = uSystolicPE_413_io_mac_done_d;
    mac_done_x_11[11] = uSystolicPE_414_io_mac_done_d;
    mac_done_x_11[12] = uSystolicPE_415_io_mac_done_d;
    mac_done_x_11[13] = uSystolicPE_416_io_mac_done_d;
    mac_done_x_11[14] = uSystolicPE_417_io_mac_done_d;
    mac_done_x_11[15] = uSystolicPE_418_io_mac_done_d;
    mac_done_x_11[16] = uSystolicPE_419_io_mac_done_d;
  end

  always @(*) begin
    enable_w_x_11[0] = io_enable_w[11];
    enable_w_x_11[1] = uSystolicPE_250_io_enable_w_d;
    enable_w_x_11[2] = uSystolicPE_265_io_enable_w_d;
    enable_w_x_11[3] = uSystolicPE_280_io_enable_w_d;
    enable_w_x_11[4] = uSystolicPE_295_io_enable_w_d;
    enable_w_x_11[5] = uSystolicPE_310_io_enable_w_d;
    enable_w_x_11[6] = uSystolicPE_325_io_enable_w_d;
    enable_w_x_11[7] = uSystolicPE_340_io_enable_w_d;
    enable_w_x_11[8] = uSystolicPE_355_io_enable_w_d;
    enable_w_x_11[9] = uSystolicPE_370_io_enable_w_d;
    enable_w_x_11[10] = uSystolicPE_385_io_enable_w_d;
    enable_w_x_11[11] = uSystolicPE_400_io_enable_w_d;
    enable_w_x_11[12] = uSystolicPE_415_io_enable_w_d;
    enable_w_x_11[13] = uSystolicPE_430_io_enable_w_d;
    enable_w_x_11[14] = uSystolicPE_445_io_enable_w_d;
    enable_w_x_11[15] = uSystolicPE_460_io_enable_w_d;
    enable_w_x_11[16] = uSystolicPE_475_io_enable_w_d;
  end

  always @(*) begin
    clear_w_x_11[0] = io_clear_w[11];
    clear_w_x_11[1] = uSystolicPE_250_io_clear_w_d;
    clear_w_x_11[2] = uSystolicPE_265_io_clear_w_d;
    clear_w_x_11[3] = uSystolicPE_280_io_clear_w_d;
    clear_w_x_11[4] = uSystolicPE_295_io_clear_w_d;
    clear_w_x_11[5] = uSystolicPE_310_io_clear_w_d;
    clear_w_x_11[6] = uSystolicPE_325_io_clear_w_d;
    clear_w_x_11[7] = uSystolicPE_340_io_clear_w_d;
    clear_w_x_11[8] = uSystolicPE_355_io_clear_w_d;
    clear_w_x_11[9] = uSystolicPE_370_io_clear_w_d;
    clear_w_x_11[10] = uSystolicPE_385_io_clear_w_d;
    clear_w_x_11[11] = uSystolicPE_400_io_clear_w_d;
    clear_w_x_11[12] = uSystolicPE_415_io_clear_w_d;
    clear_w_x_11[13] = uSystolicPE_430_io_clear_w_d;
    clear_w_x_11[14] = uSystolicPE_445_io_clear_w_d;
    clear_w_x_11[15] = uSystolicPE_460_io_clear_w_d;
    clear_w_x_11[16] = uSystolicPE_475_io_clear_w_d;
  end

  assign wght_sign_x_11_0 = io_wght_sign[11];
  assign wght_abs_x_11_0 = io_wght_abs_11;
  always @(*) begin
    enable_o_x_11[16] = io_enable_o[11];
    enable_o_x_11[0] = uSystolicPE_250_io_enable_o_d;
    enable_o_x_11[1] = uSystolicPE_265_io_enable_o_d;
    enable_o_x_11[2] = uSystolicPE_280_io_enable_o_d;
    enable_o_x_11[3] = uSystolicPE_295_io_enable_o_d;
    enable_o_x_11[4] = uSystolicPE_310_io_enable_o_d;
    enable_o_x_11[5] = uSystolicPE_325_io_enable_o_d;
    enable_o_x_11[6] = uSystolicPE_340_io_enable_o_d;
    enable_o_x_11[7] = uSystolicPE_355_io_enable_o_d;
    enable_o_x_11[8] = uSystolicPE_370_io_enable_o_d;
    enable_o_x_11[9] = uSystolicPE_385_io_enable_o_d;
    enable_o_x_11[10] = uSystolicPE_400_io_enable_o_d;
    enable_o_x_11[11] = uSystolicPE_415_io_enable_o_d;
    enable_o_x_11[12] = uSystolicPE_430_io_enable_o_d;
    enable_o_x_11[13] = uSystolicPE_445_io_enable_o_d;
    enable_o_x_11[14] = uSystolicPE_460_io_enable_o_d;
    enable_o_x_11[15] = uSystolicPE_475_io_enable_o_d;
  end

  always @(*) begin
    clear_o_x_11[16] = io_clear_o[11];
    clear_o_x_11[0] = uSystolicPE_250_io_clear_o_d;
    clear_o_x_11[1] = uSystolicPE_265_io_clear_o_d;
    clear_o_x_11[2] = uSystolicPE_280_io_clear_o_d;
    clear_o_x_11[3] = uSystolicPE_295_io_clear_o_d;
    clear_o_x_11[4] = uSystolicPE_310_io_clear_o_d;
    clear_o_x_11[5] = uSystolicPE_325_io_clear_o_d;
    clear_o_x_11[6] = uSystolicPE_340_io_clear_o_d;
    clear_o_x_11[7] = uSystolicPE_355_io_clear_o_d;
    clear_o_x_11[8] = uSystolicPE_370_io_clear_o_d;
    clear_o_x_11[9] = uSystolicPE_385_io_clear_o_d;
    clear_o_x_11[10] = uSystolicPE_400_io_clear_o_d;
    clear_o_x_11[11] = uSystolicPE_415_io_clear_o_d;
    clear_o_x_11[12] = uSystolicPE_430_io_clear_o_d;
    clear_o_x_11[13] = uSystolicPE_445_io_clear_o_d;
    clear_o_x_11[14] = uSystolicPE_460_io_clear_o_d;
    clear_o_x_11[15] = uSystolicPE_475_io_clear_o_d;
  end

  assign io_ofm_11 = ofm_x_11_0;
  assign ofm_x_11_16 = 32'h00000000;
  always @(*) begin
    enable_i_x_12[0] = io_enable_i[12];
    enable_i_x_12[1] = uSystolicPEBorder_28_io_enable_i_d;
    enable_i_x_12[2] = uSystolicPE_420_io_enable_i_d;
    enable_i_x_12[3] = uSystolicPE_421_io_enable_i_d;
    enable_i_x_12[4] = uSystolicPE_422_io_enable_i_d;
    enable_i_x_12[5] = uSystolicPE_423_io_enable_i_d;
    enable_i_x_12[6] = uSystolicPE_424_io_enable_i_d;
    enable_i_x_12[7] = uSystolicPE_425_io_enable_i_d;
    enable_i_x_12[8] = uSystolicPE_426_io_enable_i_d;
    enable_i_x_12[9] = uSystolicPE_427_io_enable_i_d;
    enable_i_x_12[10] = uSystolicPE_428_io_enable_i_d;
    enable_i_x_12[11] = uSystolicPE_429_io_enable_i_d;
    enable_i_x_12[12] = uSystolicPE_430_io_enable_i_d;
    enable_i_x_12[13] = uSystolicPE_431_io_enable_i_d;
    enable_i_x_12[14] = uSystolicPE_432_io_enable_i_d;
    enable_i_x_12[15] = uSystolicPE_433_io_enable_i_d;
    enable_i_x_12[16] = uSystolicPE_434_io_enable_i_d;
  end

  always @(*) begin
    clear_i_x_12[0] = io_clear_i[12];
    clear_i_x_12[1] = uSystolicPEBorder_28_io_clear_i_d;
    clear_i_x_12[2] = uSystolicPE_420_io_clear_i_d;
    clear_i_x_12[3] = uSystolicPE_421_io_clear_i_d;
    clear_i_x_12[4] = uSystolicPE_422_io_clear_i_d;
    clear_i_x_12[5] = uSystolicPE_423_io_clear_i_d;
    clear_i_x_12[6] = uSystolicPE_424_io_clear_i_d;
    clear_i_x_12[7] = uSystolicPE_425_io_clear_i_d;
    clear_i_x_12[8] = uSystolicPE_426_io_clear_i_d;
    clear_i_x_12[9] = uSystolicPE_427_io_clear_i_d;
    clear_i_x_12[10] = uSystolicPE_428_io_clear_i_d;
    clear_i_x_12[11] = uSystolicPE_429_io_clear_i_d;
    clear_i_x_12[12] = uSystolicPE_430_io_clear_i_d;
    clear_i_x_12[13] = uSystolicPE_431_io_clear_i_d;
    clear_i_x_12[14] = uSystolicPE_432_io_clear_i_d;
    clear_i_x_12[15] = uSystolicPE_433_io_clear_i_d;
    clear_i_x_12[16] = uSystolicPE_434_io_clear_i_d;
  end

  always @(*) begin
    mac_done_x_12[0] = io_mac_done[12];
    mac_done_x_12[1] = uSystolicPEBorder_28_io_mac_done_d;
    mac_done_x_12[2] = uSystolicPE_420_io_mac_done_d;
    mac_done_x_12[3] = uSystolicPE_421_io_mac_done_d;
    mac_done_x_12[4] = uSystolicPE_422_io_mac_done_d;
    mac_done_x_12[5] = uSystolicPE_423_io_mac_done_d;
    mac_done_x_12[6] = uSystolicPE_424_io_mac_done_d;
    mac_done_x_12[7] = uSystolicPE_425_io_mac_done_d;
    mac_done_x_12[8] = uSystolicPE_426_io_mac_done_d;
    mac_done_x_12[9] = uSystolicPE_427_io_mac_done_d;
    mac_done_x_12[10] = uSystolicPE_428_io_mac_done_d;
    mac_done_x_12[11] = uSystolicPE_429_io_mac_done_d;
    mac_done_x_12[12] = uSystolicPE_430_io_mac_done_d;
    mac_done_x_12[13] = uSystolicPE_431_io_mac_done_d;
    mac_done_x_12[14] = uSystolicPE_432_io_mac_done_d;
    mac_done_x_12[15] = uSystolicPE_433_io_mac_done_d;
    mac_done_x_12[16] = uSystolicPE_434_io_mac_done_d;
  end

  always @(*) begin
    enable_w_x_12[0] = io_enable_w[12];
    enable_w_x_12[1] = uSystolicPE_251_io_enable_w_d;
    enable_w_x_12[2] = uSystolicPE_266_io_enable_w_d;
    enable_w_x_12[3] = uSystolicPE_281_io_enable_w_d;
    enable_w_x_12[4] = uSystolicPE_296_io_enable_w_d;
    enable_w_x_12[5] = uSystolicPE_311_io_enable_w_d;
    enable_w_x_12[6] = uSystolicPE_326_io_enable_w_d;
    enable_w_x_12[7] = uSystolicPE_341_io_enable_w_d;
    enable_w_x_12[8] = uSystolicPE_356_io_enable_w_d;
    enable_w_x_12[9] = uSystolicPE_371_io_enable_w_d;
    enable_w_x_12[10] = uSystolicPE_386_io_enable_w_d;
    enable_w_x_12[11] = uSystolicPE_401_io_enable_w_d;
    enable_w_x_12[12] = uSystolicPE_416_io_enable_w_d;
    enable_w_x_12[13] = uSystolicPE_431_io_enable_w_d;
    enable_w_x_12[14] = uSystolicPE_446_io_enable_w_d;
    enable_w_x_12[15] = uSystolicPE_461_io_enable_w_d;
    enable_w_x_12[16] = uSystolicPE_476_io_enable_w_d;
  end

  always @(*) begin
    clear_w_x_12[0] = io_clear_w[12];
    clear_w_x_12[1] = uSystolicPE_251_io_clear_w_d;
    clear_w_x_12[2] = uSystolicPE_266_io_clear_w_d;
    clear_w_x_12[3] = uSystolicPE_281_io_clear_w_d;
    clear_w_x_12[4] = uSystolicPE_296_io_clear_w_d;
    clear_w_x_12[5] = uSystolicPE_311_io_clear_w_d;
    clear_w_x_12[6] = uSystolicPE_326_io_clear_w_d;
    clear_w_x_12[7] = uSystolicPE_341_io_clear_w_d;
    clear_w_x_12[8] = uSystolicPE_356_io_clear_w_d;
    clear_w_x_12[9] = uSystolicPE_371_io_clear_w_d;
    clear_w_x_12[10] = uSystolicPE_386_io_clear_w_d;
    clear_w_x_12[11] = uSystolicPE_401_io_clear_w_d;
    clear_w_x_12[12] = uSystolicPE_416_io_clear_w_d;
    clear_w_x_12[13] = uSystolicPE_431_io_clear_w_d;
    clear_w_x_12[14] = uSystolicPE_446_io_clear_w_d;
    clear_w_x_12[15] = uSystolicPE_461_io_clear_w_d;
    clear_w_x_12[16] = uSystolicPE_476_io_clear_w_d;
  end

  assign wght_sign_x_12_0 = io_wght_sign[12];
  assign wght_abs_x_12_0 = io_wght_abs_12;
  always @(*) begin
    enable_o_x_12[16] = io_enable_o[12];
    enable_o_x_12[0] = uSystolicPE_251_io_enable_o_d;
    enable_o_x_12[1] = uSystolicPE_266_io_enable_o_d;
    enable_o_x_12[2] = uSystolicPE_281_io_enable_o_d;
    enable_o_x_12[3] = uSystolicPE_296_io_enable_o_d;
    enable_o_x_12[4] = uSystolicPE_311_io_enable_o_d;
    enable_o_x_12[5] = uSystolicPE_326_io_enable_o_d;
    enable_o_x_12[6] = uSystolicPE_341_io_enable_o_d;
    enable_o_x_12[7] = uSystolicPE_356_io_enable_o_d;
    enable_o_x_12[8] = uSystolicPE_371_io_enable_o_d;
    enable_o_x_12[9] = uSystolicPE_386_io_enable_o_d;
    enable_o_x_12[10] = uSystolicPE_401_io_enable_o_d;
    enable_o_x_12[11] = uSystolicPE_416_io_enable_o_d;
    enable_o_x_12[12] = uSystolicPE_431_io_enable_o_d;
    enable_o_x_12[13] = uSystolicPE_446_io_enable_o_d;
    enable_o_x_12[14] = uSystolicPE_461_io_enable_o_d;
    enable_o_x_12[15] = uSystolicPE_476_io_enable_o_d;
  end

  always @(*) begin
    clear_o_x_12[16] = io_clear_o[12];
    clear_o_x_12[0] = uSystolicPE_251_io_clear_o_d;
    clear_o_x_12[1] = uSystolicPE_266_io_clear_o_d;
    clear_o_x_12[2] = uSystolicPE_281_io_clear_o_d;
    clear_o_x_12[3] = uSystolicPE_296_io_clear_o_d;
    clear_o_x_12[4] = uSystolicPE_311_io_clear_o_d;
    clear_o_x_12[5] = uSystolicPE_326_io_clear_o_d;
    clear_o_x_12[6] = uSystolicPE_341_io_clear_o_d;
    clear_o_x_12[7] = uSystolicPE_356_io_clear_o_d;
    clear_o_x_12[8] = uSystolicPE_371_io_clear_o_d;
    clear_o_x_12[9] = uSystolicPE_386_io_clear_o_d;
    clear_o_x_12[10] = uSystolicPE_401_io_clear_o_d;
    clear_o_x_12[11] = uSystolicPE_416_io_clear_o_d;
    clear_o_x_12[12] = uSystolicPE_431_io_clear_o_d;
    clear_o_x_12[13] = uSystolicPE_446_io_clear_o_d;
    clear_o_x_12[14] = uSystolicPE_461_io_clear_o_d;
    clear_o_x_12[15] = uSystolicPE_476_io_clear_o_d;
  end

  assign io_ofm_12 = ofm_x_12_0;
  assign ofm_x_12_16 = 32'h00000000;
  always @(*) begin
    enable_i_x_13[0] = io_enable_i[13];
    enable_i_x_13[1] = uSystolicPEBorder_29_io_enable_i_d;
    enable_i_x_13[2] = uSystolicPE_435_io_enable_i_d;
    enable_i_x_13[3] = uSystolicPE_436_io_enable_i_d;
    enable_i_x_13[4] = uSystolicPE_437_io_enable_i_d;
    enable_i_x_13[5] = uSystolicPE_438_io_enable_i_d;
    enable_i_x_13[6] = uSystolicPE_439_io_enable_i_d;
    enable_i_x_13[7] = uSystolicPE_440_io_enable_i_d;
    enable_i_x_13[8] = uSystolicPE_441_io_enable_i_d;
    enable_i_x_13[9] = uSystolicPE_442_io_enable_i_d;
    enable_i_x_13[10] = uSystolicPE_443_io_enable_i_d;
    enable_i_x_13[11] = uSystolicPE_444_io_enable_i_d;
    enable_i_x_13[12] = uSystolicPE_445_io_enable_i_d;
    enable_i_x_13[13] = uSystolicPE_446_io_enable_i_d;
    enable_i_x_13[14] = uSystolicPE_447_io_enable_i_d;
    enable_i_x_13[15] = uSystolicPE_448_io_enable_i_d;
    enable_i_x_13[16] = uSystolicPE_449_io_enable_i_d;
  end

  always @(*) begin
    clear_i_x_13[0] = io_clear_i[13];
    clear_i_x_13[1] = uSystolicPEBorder_29_io_clear_i_d;
    clear_i_x_13[2] = uSystolicPE_435_io_clear_i_d;
    clear_i_x_13[3] = uSystolicPE_436_io_clear_i_d;
    clear_i_x_13[4] = uSystolicPE_437_io_clear_i_d;
    clear_i_x_13[5] = uSystolicPE_438_io_clear_i_d;
    clear_i_x_13[6] = uSystolicPE_439_io_clear_i_d;
    clear_i_x_13[7] = uSystolicPE_440_io_clear_i_d;
    clear_i_x_13[8] = uSystolicPE_441_io_clear_i_d;
    clear_i_x_13[9] = uSystolicPE_442_io_clear_i_d;
    clear_i_x_13[10] = uSystolicPE_443_io_clear_i_d;
    clear_i_x_13[11] = uSystolicPE_444_io_clear_i_d;
    clear_i_x_13[12] = uSystolicPE_445_io_clear_i_d;
    clear_i_x_13[13] = uSystolicPE_446_io_clear_i_d;
    clear_i_x_13[14] = uSystolicPE_447_io_clear_i_d;
    clear_i_x_13[15] = uSystolicPE_448_io_clear_i_d;
    clear_i_x_13[16] = uSystolicPE_449_io_clear_i_d;
  end

  always @(*) begin
    mac_done_x_13[0] = io_mac_done[13];
    mac_done_x_13[1] = uSystolicPEBorder_29_io_mac_done_d;
    mac_done_x_13[2] = uSystolicPE_435_io_mac_done_d;
    mac_done_x_13[3] = uSystolicPE_436_io_mac_done_d;
    mac_done_x_13[4] = uSystolicPE_437_io_mac_done_d;
    mac_done_x_13[5] = uSystolicPE_438_io_mac_done_d;
    mac_done_x_13[6] = uSystolicPE_439_io_mac_done_d;
    mac_done_x_13[7] = uSystolicPE_440_io_mac_done_d;
    mac_done_x_13[8] = uSystolicPE_441_io_mac_done_d;
    mac_done_x_13[9] = uSystolicPE_442_io_mac_done_d;
    mac_done_x_13[10] = uSystolicPE_443_io_mac_done_d;
    mac_done_x_13[11] = uSystolicPE_444_io_mac_done_d;
    mac_done_x_13[12] = uSystolicPE_445_io_mac_done_d;
    mac_done_x_13[13] = uSystolicPE_446_io_mac_done_d;
    mac_done_x_13[14] = uSystolicPE_447_io_mac_done_d;
    mac_done_x_13[15] = uSystolicPE_448_io_mac_done_d;
    mac_done_x_13[16] = uSystolicPE_449_io_mac_done_d;
  end

  always @(*) begin
    enable_w_x_13[0] = io_enable_w[13];
    enable_w_x_13[1] = uSystolicPE_252_io_enable_w_d;
    enable_w_x_13[2] = uSystolicPE_267_io_enable_w_d;
    enable_w_x_13[3] = uSystolicPE_282_io_enable_w_d;
    enable_w_x_13[4] = uSystolicPE_297_io_enable_w_d;
    enable_w_x_13[5] = uSystolicPE_312_io_enable_w_d;
    enable_w_x_13[6] = uSystolicPE_327_io_enable_w_d;
    enable_w_x_13[7] = uSystolicPE_342_io_enable_w_d;
    enable_w_x_13[8] = uSystolicPE_357_io_enable_w_d;
    enable_w_x_13[9] = uSystolicPE_372_io_enable_w_d;
    enable_w_x_13[10] = uSystolicPE_387_io_enable_w_d;
    enable_w_x_13[11] = uSystolicPE_402_io_enable_w_d;
    enable_w_x_13[12] = uSystolicPE_417_io_enable_w_d;
    enable_w_x_13[13] = uSystolicPE_432_io_enable_w_d;
    enable_w_x_13[14] = uSystolicPE_447_io_enable_w_d;
    enable_w_x_13[15] = uSystolicPE_462_io_enable_w_d;
    enable_w_x_13[16] = uSystolicPE_477_io_enable_w_d;
  end

  always @(*) begin
    clear_w_x_13[0] = io_clear_w[13];
    clear_w_x_13[1] = uSystolicPE_252_io_clear_w_d;
    clear_w_x_13[2] = uSystolicPE_267_io_clear_w_d;
    clear_w_x_13[3] = uSystolicPE_282_io_clear_w_d;
    clear_w_x_13[4] = uSystolicPE_297_io_clear_w_d;
    clear_w_x_13[5] = uSystolicPE_312_io_clear_w_d;
    clear_w_x_13[6] = uSystolicPE_327_io_clear_w_d;
    clear_w_x_13[7] = uSystolicPE_342_io_clear_w_d;
    clear_w_x_13[8] = uSystolicPE_357_io_clear_w_d;
    clear_w_x_13[9] = uSystolicPE_372_io_clear_w_d;
    clear_w_x_13[10] = uSystolicPE_387_io_clear_w_d;
    clear_w_x_13[11] = uSystolicPE_402_io_clear_w_d;
    clear_w_x_13[12] = uSystolicPE_417_io_clear_w_d;
    clear_w_x_13[13] = uSystolicPE_432_io_clear_w_d;
    clear_w_x_13[14] = uSystolicPE_447_io_clear_w_d;
    clear_w_x_13[15] = uSystolicPE_462_io_clear_w_d;
    clear_w_x_13[16] = uSystolicPE_477_io_clear_w_d;
  end

  assign wght_sign_x_13_0 = io_wght_sign[13];
  assign wght_abs_x_13_0 = io_wght_abs_13;
  always @(*) begin
    enable_o_x_13[16] = io_enable_o[13];
    enable_o_x_13[0] = uSystolicPE_252_io_enable_o_d;
    enable_o_x_13[1] = uSystolicPE_267_io_enable_o_d;
    enable_o_x_13[2] = uSystolicPE_282_io_enable_o_d;
    enable_o_x_13[3] = uSystolicPE_297_io_enable_o_d;
    enable_o_x_13[4] = uSystolicPE_312_io_enable_o_d;
    enable_o_x_13[5] = uSystolicPE_327_io_enable_o_d;
    enable_o_x_13[6] = uSystolicPE_342_io_enable_o_d;
    enable_o_x_13[7] = uSystolicPE_357_io_enable_o_d;
    enable_o_x_13[8] = uSystolicPE_372_io_enable_o_d;
    enable_o_x_13[9] = uSystolicPE_387_io_enable_o_d;
    enable_o_x_13[10] = uSystolicPE_402_io_enable_o_d;
    enable_o_x_13[11] = uSystolicPE_417_io_enable_o_d;
    enable_o_x_13[12] = uSystolicPE_432_io_enable_o_d;
    enable_o_x_13[13] = uSystolicPE_447_io_enable_o_d;
    enable_o_x_13[14] = uSystolicPE_462_io_enable_o_d;
    enable_o_x_13[15] = uSystolicPE_477_io_enable_o_d;
  end

  always @(*) begin
    clear_o_x_13[16] = io_clear_o[13];
    clear_o_x_13[0] = uSystolicPE_252_io_clear_o_d;
    clear_o_x_13[1] = uSystolicPE_267_io_clear_o_d;
    clear_o_x_13[2] = uSystolicPE_282_io_clear_o_d;
    clear_o_x_13[3] = uSystolicPE_297_io_clear_o_d;
    clear_o_x_13[4] = uSystolicPE_312_io_clear_o_d;
    clear_o_x_13[5] = uSystolicPE_327_io_clear_o_d;
    clear_o_x_13[6] = uSystolicPE_342_io_clear_o_d;
    clear_o_x_13[7] = uSystolicPE_357_io_clear_o_d;
    clear_o_x_13[8] = uSystolicPE_372_io_clear_o_d;
    clear_o_x_13[9] = uSystolicPE_387_io_clear_o_d;
    clear_o_x_13[10] = uSystolicPE_402_io_clear_o_d;
    clear_o_x_13[11] = uSystolicPE_417_io_clear_o_d;
    clear_o_x_13[12] = uSystolicPE_432_io_clear_o_d;
    clear_o_x_13[13] = uSystolicPE_447_io_clear_o_d;
    clear_o_x_13[14] = uSystolicPE_462_io_clear_o_d;
    clear_o_x_13[15] = uSystolicPE_477_io_clear_o_d;
  end

  assign io_ofm_13 = ofm_x_13_0;
  assign ofm_x_13_16 = 32'h00000000;
  always @(*) begin
    enable_i_x_14[0] = io_enable_i[14];
    enable_i_x_14[1] = uSystolicPEBorder_30_io_enable_i_d;
    enable_i_x_14[2] = uSystolicPE_450_io_enable_i_d;
    enable_i_x_14[3] = uSystolicPE_451_io_enable_i_d;
    enable_i_x_14[4] = uSystolicPE_452_io_enable_i_d;
    enable_i_x_14[5] = uSystolicPE_453_io_enable_i_d;
    enable_i_x_14[6] = uSystolicPE_454_io_enable_i_d;
    enable_i_x_14[7] = uSystolicPE_455_io_enable_i_d;
    enable_i_x_14[8] = uSystolicPE_456_io_enable_i_d;
    enable_i_x_14[9] = uSystolicPE_457_io_enable_i_d;
    enable_i_x_14[10] = uSystolicPE_458_io_enable_i_d;
    enable_i_x_14[11] = uSystolicPE_459_io_enable_i_d;
    enable_i_x_14[12] = uSystolicPE_460_io_enable_i_d;
    enable_i_x_14[13] = uSystolicPE_461_io_enable_i_d;
    enable_i_x_14[14] = uSystolicPE_462_io_enable_i_d;
    enable_i_x_14[15] = uSystolicPE_463_io_enable_i_d;
    enable_i_x_14[16] = uSystolicPE_464_io_enable_i_d;
  end

  always @(*) begin
    clear_i_x_14[0] = io_clear_i[14];
    clear_i_x_14[1] = uSystolicPEBorder_30_io_clear_i_d;
    clear_i_x_14[2] = uSystolicPE_450_io_clear_i_d;
    clear_i_x_14[3] = uSystolicPE_451_io_clear_i_d;
    clear_i_x_14[4] = uSystolicPE_452_io_clear_i_d;
    clear_i_x_14[5] = uSystolicPE_453_io_clear_i_d;
    clear_i_x_14[6] = uSystolicPE_454_io_clear_i_d;
    clear_i_x_14[7] = uSystolicPE_455_io_clear_i_d;
    clear_i_x_14[8] = uSystolicPE_456_io_clear_i_d;
    clear_i_x_14[9] = uSystolicPE_457_io_clear_i_d;
    clear_i_x_14[10] = uSystolicPE_458_io_clear_i_d;
    clear_i_x_14[11] = uSystolicPE_459_io_clear_i_d;
    clear_i_x_14[12] = uSystolicPE_460_io_clear_i_d;
    clear_i_x_14[13] = uSystolicPE_461_io_clear_i_d;
    clear_i_x_14[14] = uSystolicPE_462_io_clear_i_d;
    clear_i_x_14[15] = uSystolicPE_463_io_clear_i_d;
    clear_i_x_14[16] = uSystolicPE_464_io_clear_i_d;
  end

  always @(*) begin
    mac_done_x_14[0] = io_mac_done[14];
    mac_done_x_14[1] = uSystolicPEBorder_30_io_mac_done_d;
    mac_done_x_14[2] = uSystolicPE_450_io_mac_done_d;
    mac_done_x_14[3] = uSystolicPE_451_io_mac_done_d;
    mac_done_x_14[4] = uSystolicPE_452_io_mac_done_d;
    mac_done_x_14[5] = uSystolicPE_453_io_mac_done_d;
    mac_done_x_14[6] = uSystolicPE_454_io_mac_done_d;
    mac_done_x_14[7] = uSystolicPE_455_io_mac_done_d;
    mac_done_x_14[8] = uSystolicPE_456_io_mac_done_d;
    mac_done_x_14[9] = uSystolicPE_457_io_mac_done_d;
    mac_done_x_14[10] = uSystolicPE_458_io_mac_done_d;
    mac_done_x_14[11] = uSystolicPE_459_io_mac_done_d;
    mac_done_x_14[12] = uSystolicPE_460_io_mac_done_d;
    mac_done_x_14[13] = uSystolicPE_461_io_mac_done_d;
    mac_done_x_14[14] = uSystolicPE_462_io_mac_done_d;
    mac_done_x_14[15] = uSystolicPE_463_io_mac_done_d;
    mac_done_x_14[16] = uSystolicPE_464_io_mac_done_d;
  end

  always @(*) begin
    enable_w_x_14[0] = io_enable_w[14];
    enable_w_x_14[1] = uSystolicPE_253_io_enable_w_d;
    enable_w_x_14[2] = uSystolicPE_268_io_enable_w_d;
    enable_w_x_14[3] = uSystolicPE_283_io_enable_w_d;
    enable_w_x_14[4] = uSystolicPE_298_io_enable_w_d;
    enable_w_x_14[5] = uSystolicPE_313_io_enable_w_d;
    enable_w_x_14[6] = uSystolicPE_328_io_enable_w_d;
    enable_w_x_14[7] = uSystolicPE_343_io_enable_w_d;
    enable_w_x_14[8] = uSystolicPE_358_io_enable_w_d;
    enable_w_x_14[9] = uSystolicPE_373_io_enable_w_d;
    enable_w_x_14[10] = uSystolicPE_388_io_enable_w_d;
    enable_w_x_14[11] = uSystolicPE_403_io_enable_w_d;
    enable_w_x_14[12] = uSystolicPE_418_io_enable_w_d;
    enable_w_x_14[13] = uSystolicPE_433_io_enable_w_d;
    enable_w_x_14[14] = uSystolicPE_448_io_enable_w_d;
    enable_w_x_14[15] = uSystolicPE_463_io_enable_w_d;
    enable_w_x_14[16] = uSystolicPE_478_io_enable_w_d;
  end

  always @(*) begin
    clear_w_x_14[0] = io_clear_w[14];
    clear_w_x_14[1] = uSystolicPE_253_io_clear_w_d;
    clear_w_x_14[2] = uSystolicPE_268_io_clear_w_d;
    clear_w_x_14[3] = uSystolicPE_283_io_clear_w_d;
    clear_w_x_14[4] = uSystolicPE_298_io_clear_w_d;
    clear_w_x_14[5] = uSystolicPE_313_io_clear_w_d;
    clear_w_x_14[6] = uSystolicPE_328_io_clear_w_d;
    clear_w_x_14[7] = uSystolicPE_343_io_clear_w_d;
    clear_w_x_14[8] = uSystolicPE_358_io_clear_w_d;
    clear_w_x_14[9] = uSystolicPE_373_io_clear_w_d;
    clear_w_x_14[10] = uSystolicPE_388_io_clear_w_d;
    clear_w_x_14[11] = uSystolicPE_403_io_clear_w_d;
    clear_w_x_14[12] = uSystolicPE_418_io_clear_w_d;
    clear_w_x_14[13] = uSystolicPE_433_io_clear_w_d;
    clear_w_x_14[14] = uSystolicPE_448_io_clear_w_d;
    clear_w_x_14[15] = uSystolicPE_463_io_clear_w_d;
    clear_w_x_14[16] = uSystolicPE_478_io_clear_w_d;
  end

  assign wght_sign_x_14_0 = io_wght_sign[14];
  assign wght_abs_x_14_0 = io_wght_abs_14;
  always @(*) begin
    enable_o_x_14[16] = io_enable_o[14];
    enable_o_x_14[0] = uSystolicPE_253_io_enable_o_d;
    enable_o_x_14[1] = uSystolicPE_268_io_enable_o_d;
    enable_o_x_14[2] = uSystolicPE_283_io_enable_o_d;
    enable_o_x_14[3] = uSystolicPE_298_io_enable_o_d;
    enable_o_x_14[4] = uSystolicPE_313_io_enable_o_d;
    enable_o_x_14[5] = uSystolicPE_328_io_enable_o_d;
    enable_o_x_14[6] = uSystolicPE_343_io_enable_o_d;
    enable_o_x_14[7] = uSystolicPE_358_io_enable_o_d;
    enable_o_x_14[8] = uSystolicPE_373_io_enable_o_d;
    enable_o_x_14[9] = uSystolicPE_388_io_enable_o_d;
    enable_o_x_14[10] = uSystolicPE_403_io_enable_o_d;
    enable_o_x_14[11] = uSystolicPE_418_io_enable_o_d;
    enable_o_x_14[12] = uSystolicPE_433_io_enable_o_d;
    enable_o_x_14[13] = uSystolicPE_448_io_enable_o_d;
    enable_o_x_14[14] = uSystolicPE_463_io_enable_o_d;
    enable_o_x_14[15] = uSystolicPE_478_io_enable_o_d;
  end

  always @(*) begin
    clear_o_x_14[16] = io_clear_o[14];
    clear_o_x_14[0] = uSystolicPE_253_io_clear_o_d;
    clear_o_x_14[1] = uSystolicPE_268_io_clear_o_d;
    clear_o_x_14[2] = uSystolicPE_283_io_clear_o_d;
    clear_o_x_14[3] = uSystolicPE_298_io_clear_o_d;
    clear_o_x_14[4] = uSystolicPE_313_io_clear_o_d;
    clear_o_x_14[5] = uSystolicPE_328_io_clear_o_d;
    clear_o_x_14[6] = uSystolicPE_343_io_clear_o_d;
    clear_o_x_14[7] = uSystolicPE_358_io_clear_o_d;
    clear_o_x_14[8] = uSystolicPE_373_io_clear_o_d;
    clear_o_x_14[9] = uSystolicPE_388_io_clear_o_d;
    clear_o_x_14[10] = uSystolicPE_403_io_clear_o_d;
    clear_o_x_14[11] = uSystolicPE_418_io_clear_o_d;
    clear_o_x_14[12] = uSystolicPE_433_io_clear_o_d;
    clear_o_x_14[13] = uSystolicPE_448_io_clear_o_d;
    clear_o_x_14[14] = uSystolicPE_463_io_clear_o_d;
    clear_o_x_14[15] = uSystolicPE_478_io_clear_o_d;
  end

  assign io_ofm_14 = ofm_x_14_0;
  assign ofm_x_14_16 = 32'h00000000;
  always @(*) begin
    enable_i_x_15[0] = io_enable_i[15];
    enable_i_x_15[1] = uSystolicPEBorder_31_io_enable_i_d;
    enable_i_x_15[2] = uSystolicPE_465_io_enable_i_d;
    enable_i_x_15[3] = uSystolicPE_466_io_enable_i_d;
    enable_i_x_15[4] = uSystolicPE_467_io_enable_i_d;
    enable_i_x_15[5] = uSystolicPE_468_io_enable_i_d;
    enable_i_x_15[6] = uSystolicPE_469_io_enable_i_d;
    enable_i_x_15[7] = uSystolicPE_470_io_enable_i_d;
    enable_i_x_15[8] = uSystolicPE_471_io_enable_i_d;
    enable_i_x_15[9] = uSystolicPE_472_io_enable_i_d;
    enable_i_x_15[10] = uSystolicPE_473_io_enable_i_d;
    enable_i_x_15[11] = uSystolicPE_474_io_enable_i_d;
    enable_i_x_15[12] = uSystolicPE_475_io_enable_i_d;
    enable_i_x_15[13] = uSystolicPE_476_io_enable_i_d;
    enable_i_x_15[14] = uSystolicPE_477_io_enable_i_d;
    enable_i_x_15[15] = uSystolicPE_478_io_enable_i_d;
    enable_i_x_15[16] = uSystolicPE_479_io_enable_i_d;
  end

  always @(*) begin
    clear_i_x_15[0] = io_clear_i[15];
    clear_i_x_15[1] = uSystolicPEBorder_31_io_clear_i_d;
    clear_i_x_15[2] = uSystolicPE_465_io_clear_i_d;
    clear_i_x_15[3] = uSystolicPE_466_io_clear_i_d;
    clear_i_x_15[4] = uSystolicPE_467_io_clear_i_d;
    clear_i_x_15[5] = uSystolicPE_468_io_clear_i_d;
    clear_i_x_15[6] = uSystolicPE_469_io_clear_i_d;
    clear_i_x_15[7] = uSystolicPE_470_io_clear_i_d;
    clear_i_x_15[8] = uSystolicPE_471_io_clear_i_d;
    clear_i_x_15[9] = uSystolicPE_472_io_clear_i_d;
    clear_i_x_15[10] = uSystolicPE_473_io_clear_i_d;
    clear_i_x_15[11] = uSystolicPE_474_io_clear_i_d;
    clear_i_x_15[12] = uSystolicPE_475_io_clear_i_d;
    clear_i_x_15[13] = uSystolicPE_476_io_clear_i_d;
    clear_i_x_15[14] = uSystolicPE_477_io_clear_i_d;
    clear_i_x_15[15] = uSystolicPE_478_io_clear_i_d;
    clear_i_x_15[16] = uSystolicPE_479_io_clear_i_d;
  end

  always @(*) begin
    mac_done_x_15[0] = io_mac_done[15];
    mac_done_x_15[1] = uSystolicPEBorder_31_io_mac_done_d;
    mac_done_x_15[2] = uSystolicPE_465_io_mac_done_d;
    mac_done_x_15[3] = uSystolicPE_466_io_mac_done_d;
    mac_done_x_15[4] = uSystolicPE_467_io_mac_done_d;
    mac_done_x_15[5] = uSystolicPE_468_io_mac_done_d;
    mac_done_x_15[6] = uSystolicPE_469_io_mac_done_d;
    mac_done_x_15[7] = uSystolicPE_470_io_mac_done_d;
    mac_done_x_15[8] = uSystolicPE_471_io_mac_done_d;
    mac_done_x_15[9] = uSystolicPE_472_io_mac_done_d;
    mac_done_x_15[10] = uSystolicPE_473_io_mac_done_d;
    mac_done_x_15[11] = uSystolicPE_474_io_mac_done_d;
    mac_done_x_15[12] = uSystolicPE_475_io_mac_done_d;
    mac_done_x_15[13] = uSystolicPE_476_io_mac_done_d;
    mac_done_x_15[14] = uSystolicPE_477_io_mac_done_d;
    mac_done_x_15[15] = uSystolicPE_478_io_mac_done_d;
    mac_done_x_15[16] = uSystolicPE_479_io_mac_done_d;
  end

  always @(*) begin
    enable_w_x_15[0] = io_enable_w[15];
    enable_w_x_15[1] = uSystolicPE_254_io_enable_w_d;
    enable_w_x_15[2] = uSystolicPE_269_io_enable_w_d;
    enable_w_x_15[3] = uSystolicPE_284_io_enable_w_d;
    enable_w_x_15[4] = uSystolicPE_299_io_enable_w_d;
    enable_w_x_15[5] = uSystolicPE_314_io_enable_w_d;
    enable_w_x_15[6] = uSystolicPE_329_io_enable_w_d;
    enable_w_x_15[7] = uSystolicPE_344_io_enable_w_d;
    enable_w_x_15[8] = uSystolicPE_359_io_enable_w_d;
    enable_w_x_15[9] = uSystolicPE_374_io_enable_w_d;
    enable_w_x_15[10] = uSystolicPE_389_io_enable_w_d;
    enable_w_x_15[11] = uSystolicPE_404_io_enable_w_d;
    enable_w_x_15[12] = uSystolicPE_419_io_enable_w_d;
    enable_w_x_15[13] = uSystolicPE_434_io_enable_w_d;
    enable_w_x_15[14] = uSystolicPE_449_io_enable_w_d;
    enable_w_x_15[15] = uSystolicPE_464_io_enable_w_d;
    enable_w_x_15[16] = uSystolicPE_479_io_enable_w_d;
  end

  always @(*) begin
    clear_w_x_15[0] = io_clear_w[15];
    clear_w_x_15[1] = uSystolicPE_254_io_clear_w_d;
    clear_w_x_15[2] = uSystolicPE_269_io_clear_w_d;
    clear_w_x_15[3] = uSystolicPE_284_io_clear_w_d;
    clear_w_x_15[4] = uSystolicPE_299_io_clear_w_d;
    clear_w_x_15[5] = uSystolicPE_314_io_clear_w_d;
    clear_w_x_15[6] = uSystolicPE_329_io_clear_w_d;
    clear_w_x_15[7] = uSystolicPE_344_io_clear_w_d;
    clear_w_x_15[8] = uSystolicPE_359_io_clear_w_d;
    clear_w_x_15[9] = uSystolicPE_374_io_clear_w_d;
    clear_w_x_15[10] = uSystolicPE_389_io_clear_w_d;
    clear_w_x_15[11] = uSystolicPE_404_io_clear_w_d;
    clear_w_x_15[12] = uSystolicPE_419_io_clear_w_d;
    clear_w_x_15[13] = uSystolicPE_434_io_clear_w_d;
    clear_w_x_15[14] = uSystolicPE_449_io_clear_w_d;
    clear_w_x_15[15] = uSystolicPE_464_io_clear_w_d;
    clear_w_x_15[16] = uSystolicPE_479_io_clear_w_d;
  end

  assign wght_sign_x_15_0 = io_wght_sign[15];
  assign wght_abs_x_15_0 = io_wght_abs_15;
  always @(*) begin
    enable_o_x_15[16] = io_enable_o[15];
    enable_o_x_15[0] = uSystolicPE_254_io_enable_o_d;
    enable_o_x_15[1] = uSystolicPE_269_io_enable_o_d;
    enable_o_x_15[2] = uSystolicPE_284_io_enable_o_d;
    enable_o_x_15[3] = uSystolicPE_299_io_enable_o_d;
    enable_o_x_15[4] = uSystolicPE_314_io_enable_o_d;
    enable_o_x_15[5] = uSystolicPE_329_io_enable_o_d;
    enable_o_x_15[6] = uSystolicPE_344_io_enable_o_d;
    enable_o_x_15[7] = uSystolicPE_359_io_enable_o_d;
    enable_o_x_15[8] = uSystolicPE_374_io_enable_o_d;
    enable_o_x_15[9] = uSystolicPE_389_io_enable_o_d;
    enable_o_x_15[10] = uSystolicPE_404_io_enable_o_d;
    enable_o_x_15[11] = uSystolicPE_419_io_enable_o_d;
    enable_o_x_15[12] = uSystolicPE_434_io_enable_o_d;
    enable_o_x_15[13] = uSystolicPE_449_io_enable_o_d;
    enable_o_x_15[14] = uSystolicPE_464_io_enable_o_d;
    enable_o_x_15[15] = uSystolicPE_479_io_enable_o_d;
  end

  always @(*) begin
    clear_o_x_15[16] = io_clear_o[15];
    clear_o_x_15[0] = uSystolicPE_254_io_clear_o_d;
    clear_o_x_15[1] = uSystolicPE_269_io_clear_o_d;
    clear_o_x_15[2] = uSystolicPE_284_io_clear_o_d;
    clear_o_x_15[3] = uSystolicPE_299_io_clear_o_d;
    clear_o_x_15[4] = uSystolicPE_314_io_clear_o_d;
    clear_o_x_15[5] = uSystolicPE_329_io_clear_o_d;
    clear_o_x_15[6] = uSystolicPE_344_io_clear_o_d;
    clear_o_x_15[7] = uSystolicPE_359_io_clear_o_d;
    clear_o_x_15[8] = uSystolicPE_374_io_clear_o_d;
    clear_o_x_15[9] = uSystolicPE_389_io_clear_o_d;
    clear_o_x_15[10] = uSystolicPE_404_io_clear_o_d;
    clear_o_x_15[11] = uSystolicPE_419_io_clear_o_d;
    clear_o_x_15[12] = uSystolicPE_434_io_clear_o_d;
    clear_o_x_15[13] = uSystolicPE_449_io_clear_o_d;
    clear_o_x_15[14] = uSystolicPE_464_io_clear_o_d;
    clear_o_x_15[15] = uSystolicPE_479_io_clear_o_d;
  end

  assign io_ofm_15 = ofm_x_15_0;
  assign ofm_x_15_16 = 32'h00000000;
  assign uSystolicPEBorder_16_io_mac_done = mac_done_x_0[0];
  assign uSystolicPEBorder_16_io_enable_i = enable_i_x_0[0];
  assign uSystolicPEBorder_16_io_clear_i = clear_i_x_0[0];
  assign ifm_sign_x_0_1 = uSystolicPEBorder_16_io_ifm_sign_d;
  assign ifm_dff_x_0_1 = uSystolicPEBorder_16_io_ifm_dff_d;
  assign uSystolicPEBorder_16_io_enable_w = enable_w_x_0[0];
  assign uSystolicPEBorder_16_io_clear_w = clear_w_x_0[0];
  assign wght_sign_x_0_1 = uSystolicPEBorder_16_io_wght_sign_d;
  assign wght_abs_x_0_1 = uSystolicPEBorder_16_io_wght_abs_d;
  assign uSystolicPEBorder_16_io_enable_o = enable_o_x_0[1];
  assign uSystolicPEBorder_16_io_clear_o = clear_o_x_0[1];
  assign ofm_x_0_0 = uSystolicPEBorder_16_io_ofm_d;
  assign randW_x_0_1 = uSystolicPEBorder_16_io_randW_d;
  assign uSystolicPE_240_io_mac_done = mac_done_x_0[1];
  assign uSystolicPE_240_io_enable_i = enable_i_x_0[1];
  assign uSystolicPE_240_io_clear_i = clear_i_x_0[1];
  assign ifm_sign_x_0_2 = uSystolicPE_240_io_ifm_sign_d;
  assign ifm_dff_x_0_2 = uSystolicPE_240_io_ifm_dff_d;
  assign uSystolicPE_240_io_enable_w = enable_w_x_1[0];
  assign uSystolicPE_240_io_clear_w = clear_w_x_1[0];
  assign wght_sign_x_1_1 = uSystolicPE_240_io_wght_sign_d;
  assign wght_abs_x_1_1 = uSystolicPE_240_io_wght_abs_d;
  assign uSystolicPE_240_io_enable_o = enable_o_x_1[1];
  assign uSystolicPE_240_io_clear_o = clear_o_x_1[1];
  assign ofm_x_1_0 = uSystolicPE_240_io_ofm_d;
  assign randW_x_0_2 = uSystolicPE_240_io_randW_d;
  assign uSystolicPE_241_io_mac_done = mac_done_x_0[2];
  assign uSystolicPE_241_io_enable_i = enable_i_x_0[2];
  assign uSystolicPE_241_io_clear_i = clear_i_x_0[2];
  assign ifm_sign_x_0_3 = uSystolicPE_241_io_ifm_sign_d;
  assign ifm_dff_x_0_3 = uSystolicPE_241_io_ifm_dff_d;
  assign uSystolicPE_241_io_enable_w = enable_w_x_2[0];
  assign uSystolicPE_241_io_clear_w = clear_w_x_2[0];
  assign wght_sign_x_2_1 = uSystolicPE_241_io_wght_sign_d;
  assign wght_abs_x_2_1 = uSystolicPE_241_io_wght_abs_d;
  assign uSystolicPE_241_io_enable_o = enable_o_x_2[1];
  assign uSystolicPE_241_io_clear_o = clear_o_x_2[1];
  assign ofm_x_2_0 = uSystolicPE_241_io_ofm_d;
  assign randW_x_0_3 = uSystolicPE_241_io_randW_d;
  assign uSystolicPE_242_io_mac_done = mac_done_x_0[3];
  assign uSystolicPE_242_io_enable_i = enable_i_x_0[3];
  assign uSystolicPE_242_io_clear_i = clear_i_x_0[3];
  assign ifm_sign_x_0_4 = uSystolicPE_242_io_ifm_sign_d;
  assign ifm_dff_x_0_4 = uSystolicPE_242_io_ifm_dff_d;
  assign uSystolicPE_242_io_enable_w = enable_w_x_3[0];
  assign uSystolicPE_242_io_clear_w = clear_w_x_3[0];
  assign wght_sign_x_3_1 = uSystolicPE_242_io_wght_sign_d;
  assign wght_abs_x_3_1 = uSystolicPE_242_io_wght_abs_d;
  assign uSystolicPE_242_io_enable_o = enable_o_x_3[1];
  assign uSystolicPE_242_io_clear_o = clear_o_x_3[1];
  assign ofm_x_3_0 = uSystolicPE_242_io_ofm_d;
  assign randW_x_0_4 = uSystolicPE_242_io_randW_d;
  assign uSystolicPE_243_io_mac_done = mac_done_x_0[4];
  assign uSystolicPE_243_io_enable_i = enable_i_x_0[4];
  assign uSystolicPE_243_io_clear_i = clear_i_x_0[4];
  assign ifm_sign_x_0_5 = uSystolicPE_243_io_ifm_sign_d;
  assign ifm_dff_x_0_5 = uSystolicPE_243_io_ifm_dff_d;
  assign uSystolicPE_243_io_enable_w = enable_w_x_4[0];
  assign uSystolicPE_243_io_clear_w = clear_w_x_4[0];
  assign wght_sign_x_4_1 = uSystolicPE_243_io_wght_sign_d;
  assign wght_abs_x_4_1 = uSystolicPE_243_io_wght_abs_d;
  assign uSystolicPE_243_io_enable_o = enable_o_x_4[1];
  assign uSystolicPE_243_io_clear_o = clear_o_x_4[1];
  assign ofm_x_4_0 = uSystolicPE_243_io_ofm_d;
  assign randW_x_0_5 = uSystolicPE_243_io_randW_d;
  assign uSystolicPE_244_io_mac_done = mac_done_x_0[5];
  assign uSystolicPE_244_io_enable_i = enable_i_x_0[5];
  assign uSystolicPE_244_io_clear_i = clear_i_x_0[5];
  assign ifm_sign_x_0_6 = uSystolicPE_244_io_ifm_sign_d;
  assign ifm_dff_x_0_6 = uSystolicPE_244_io_ifm_dff_d;
  assign uSystolicPE_244_io_enable_w = enable_w_x_5[0];
  assign uSystolicPE_244_io_clear_w = clear_w_x_5[0];
  assign wght_sign_x_5_1 = uSystolicPE_244_io_wght_sign_d;
  assign wght_abs_x_5_1 = uSystolicPE_244_io_wght_abs_d;
  assign uSystolicPE_244_io_enable_o = enable_o_x_5[1];
  assign uSystolicPE_244_io_clear_o = clear_o_x_5[1];
  assign ofm_x_5_0 = uSystolicPE_244_io_ofm_d;
  assign randW_x_0_6 = uSystolicPE_244_io_randW_d;
  assign uSystolicPE_245_io_mac_done = mac_done_x_0[6];
  assign uSystolicPE_245_io_enable_i = enable_i_x_0[6];
  assign uSystolicPE_245_io_clear_i = clear_i_x_0[6];
  assign ifm_sign_x_0_7 = uSystolicPE_245_io_ifm_sign_d;
  assign ifm_dff_x_0_7 = uSystolicPE_245_io_ifm_dff_d;
  assign uSystolicPE_245_io_enable_w = enable_w_x_6[0];
  assign uSystolicPE_245_io_clear_w = clear_w_x_6[0];
  assign wght_sign_x_6_1 = uSystolicPE_245_io_wght_sign_d;
  assign wght_abs_x_6_1 = uSystolicPE_245_io_wght_abs_d;
  assign uSystolicPE_245_io_enable_o = enable_o_x_6[1];
  assign uSystolicPE_245_io_clear_o = clear_o_x_6[1];
  assign ofm_x_6_0 = uSystolicPE_245_io_ofm_d;
  assign randW_x_0_7 = uSystolicPE_245_io_randW_d;
  assign uSystolicPE_246_io_mac_done = mac_done_x_0[7];
  assign uSystolicPE_246_io_enable_i = enable_i_x_0[7];
  assign uSystolicPE_246_io_clear_i = clear_i_x_0[7];
  assign ifm_sign_x_0_8 = uSystolicPE_246_io_ifm_sign_d;
  assign ifm_dff_x_0_8 = uSystolicPE_246_io_ifm_dff_d;
  assign uSystolicPE_246_io_enable_w = enable_w_x_7[0];
  assign uSystolicPE_246_io_clear_w = clear_w_x_7[0];
  assign wght_sign_x_7_1 = uSystolicPE_246_io_wght_sign_d;
  assign wght_abs_x_7_1 = uSystolicPE_246_io_wght_abs_d;
  assign uSystolicPE_246_io_enable_o = enable_o_x_7[1];
  assign uSystolicPE_246_io_clear_o = clear_o_x_7[1];
  assign ofm_x_7_0 = uSystolicPE_246_io_ofm_d;
  assign randW_x_0_8 = uSystolicPE_246_io_randW_d;
  assign uSystolicPE_247_io_mac_done = mac_done_x_0[8];
  assign uSystolicPE_247_io_enable_i = enable_i_x_0[8];
  assign uSystolicPE_247_io_clear_i = clear_i_x_0[8];
  assign ifm_sign_x_0_9 = uSystolicPE_247_io_ifm_sign_d;
  assign ifm_dff_x_0_9 = uSystolicPE_247_io_ifm_dff_d;
  assign uSystolicPE_247_io_enable_w = enable_w_x_8[0];
  assign uSystolicPE_247_io_clear_w = clear_w_x_8[0];
  assign wght_sign_x_8_1 = uSystolicPE_247_io_wght_sign_d;
  assign wght_abs_x_8_1 = uSystolicPE_247_io_wght_abs_d;
  assign uSystolicPE_247_io_enable_o = enable_o_x_8[1];
  assign uSystolicPE_247_io_clear_o = clear_o_x_8[1];
  assign ofm_x_8_0 = uSystolicPE_247_io_ofm_d;
  assign randW_x_0_9 = uSystolicPE_247_io_randW_d;
  assign uSystolicPE_248_io_mac_done = mac_done_x_0[9];
  assign uSystolicPE_248_io_enable_i = enable_i_x_0[9];
  assign uSystolicPE_248_io_clear_i = clear_i_x_0[9];
  assign ifm_sign_x_0_10 = uSystolicPE_248_io_ifm_sign_d;
  assign ifm_dff_x_0_10 = uSystolicPE_248_io_ifm_dff_d;
  assign uSystolicPE_248_io_enable_w = enable_w_x_9[0];
  assign uSystolicPE_248_io_clear_w = clear_w_x_9[0];
  assign wght_sign_x_9_1 = uSystolicPE_248_io_wght_sign_d;
  assign wght_abs_x_9_1 = uSystolicPE_248_io_wght_abs_d;
  assign uSystolicPE_248_io_enable_o = enable_o_x_9[1];
  assign uSystolicPE_248_io_clear_o = clear_o_x_9[1];
  assign ofm_x_9_0 = uSystolicPE_248_io_ofm_d;
  assign randW_x_0_10 = uSystolicPE_248_io_randW_d;
  assign uSystolicPE_249_io_mac_done = mac_done_x_0[10];
  assign uSystolicPE_249_io_enable_i = enable_i_x_0[10];
  assign uSystolicPE_249_io_clear_i = clear_i_x_0[10];
  assign ifm_sign_x_0_11 = uSystolicPE_249_io_ifm_sign_d;
  assign ifm_dff_x_0_11 = uSystolicPE_249_io_ifm_dff_d;
  assign uSystolicPE_249_io_enable_w = enable_w_x_10[0];
  assign uSystolicPE_249_io_clear_w = clear_w_x_10[0];
  assign wght_sign_x_10_1 = uSystolicPE_249_io_wght_sign_d;
  assign wght_abs_x_10_1 = uSystolicPE_249_io_wght_abs_d;
  assign uSystolicPE_249_io_enable_o = enable_o_x_10[1];
  assign uSystolicPE_249_io_clear_o = clear_o_x_10[1];
  assign ofm_x_10_0 = uSystolicPE_249_io_ofm_d;
  assign randW_x_0_11 = uSystolicPE_249_io_randW_d;
  assign uSystolicPE_250_io_mac_done = mac_done_x_0[11];
  assign uSystolicPE_250_io_enable_i = enable_i_x_0[11];
  assign uSystolicPE_250_io_clear_i = clear_i_x_0[11];
  assign ifm_sign_x_0_12 = uSystolicPE_250_io_ifm_sign_d;
  assign ifm_dff_x_0_12 = uSystolicPE_250_io_ifm_dff_d;
  assign uSystolicPE_250_io_enable_w = enable_w_x_11[0];
  assign uSystolicPE_250_io_clear_w = clear_w_x_11[0];
  assign wght_sign_x_11_1 = uSystolicPE_250_io_wght_sign_d;
  assign wght_abs_x_11_1 = uSystolicPE_250_io_wght_abs_d;
  assign uSystolicPE_250_io_enable_o = enable_o_x_11[1];
  assign uSystolicPE_250_io_clear_o = clear_o_x_11[1];
  assign ofm_x_11_0 = uSystolicPE_250_io_ofm_d;
  assign randW_x_0_12 = uSystolicPE_250_io_randW_d;
  assign uSystolicPE_251_io_mac_done = mac_done_x_0[12];
  assign uSystolicPE_251_io_enable_i = enable_i_x_0[12];
  assign uSystolicPE_251_io_clear_i = clear_i_x_0[12];
  assign ifm_sign_x_0_13 = uSystolicPE_251_io_ifm_sign_d;
  assign ifm_dff_x_0_13 = uSystolicPE_251_io_ifm_dff_d;
  assign uSystolicPE_251_io_enable_w = enable_w_x_12[0];
  assign uSystolicPE_251_io_clear_w = clear_w_x_12[0];
  assign wght_sign_x_12_1 = uSystolicPE_251_io_wght_sign_d;
  assign wght_abs_x_12_1 = uSystolicPE_251_io_wght_abs_d;
  assign uSystolicPE_251_io_enable_o = enable_o_x_12[1];
  assign uSystolicPE_251_io_clear_o = clear_o_x_12[1];
  assign ofm_x_12_0 = uSystolicPE_251_io_ofm_d;
  assign randW_x_0_13 = uSystolicPE_251_io_randW_d;
  assign uSystolicPE_252_io_mac_done = mac_done_x_0[13];
  assign uSystolicPE_252_io_enable_i = enable_i_x_0[13];
  assign uSystolicPE_252_io_clear_i = clear_i_x_0[13];
  assign ifm_sign_x_0_14 = uSystolicPE_252_io_ifm_sign_d;
  assign ifm_dff_x_0_14 = uSystolicPE_252_io_ifm_dff_d;
  assign uSystolicPE_252_io_enable_w = enable_w_x_13[0];
  assign uSystolicPE_252_io_clear_w = clear_w_x_13[0];
  assign wght_sign_x_13_1 = uSystolicPE_252_io_wght_sign_d;
  assign wght_abs_x_13_1 = uSystolicPE_252_io_wght_abs_d;
  assign uSystolicPE_252_io_enable_o = enable_o_x_13[1];
  assign uSystolicPE_252_io_clear_o = clear_o_x_13[1];
  assign ofm_x_13_0 = uSystolicPE_252_io_ofm_d;
  assign randW_x_0_14 = uSystolicPE_252_io_randW_d;
  assign uSystolicPE_253_io_mac_done = mac_done_x_0[14];
  assign uSystolicPE_253_io_enable_i = enable_i_x_0[14];
  assign uSystolicPE_253_io_clear_i = clear_i_x_0[14];
  assign ifm_sign_x_0_15 = uSystolicPE_253_io_ifm_sign_d;
  assign ifm_dff_x_0_15 = uSystolicPE_253_io_ifm_dff_d;
  assign uSystolicPE_253_io_enable_w = enable_w_x_14[0];
  assign uSystolicPE_253_io_clear_w = clear_w_x_14[0];
  assign wght_sign_x_14_1 = uSystolicPE_253_io_wght_sign_d;
  assign wght_abs_x_14_1 = uSystolicPE_253_io_wght_abs_d;
  assign uSystolicPE_253_io_enable_o = enable_o_x_14[1];
  assign uSystolicPE_253_io_clear_o = clear_o_x_14[1];
  assign ofm_x_14_0 = uSystolicPE_253_io_ofm_d;
  assign randW_x_0_15 = uSystolicPE_253_io_randW_d;
  assign uSystolicPE_254_io_mac_done = mac_done_x_0[15];
  assign uSystolicPE_254_io_enable_i = enable_i_x_0[15];
  assign uSystolicPE_254_io_clear_i = clear_i_x_0[15];
  assign ifm_sign_x_0_16 = uSystolicPE_254_io_ifm_sign_d;
  assign ifm_dff_x_0_16 = uSystolicPE_254_io_ifm_dff_d;
  assign uSystolicPE_254_io_enable_w = enable_w_x_15[0];
  assign uSystolicPE_254_io_clear_w = clear_w_x_15[0];
  assign wght_sign_x_15_1 = uSystolicPE_254_io_wght_sign_d;
  assign wght_abs_x_15_1 = uSystolicPE_254_io_wght_abs_d;
  assign uSystolicPE_254_io_enable_o = enable_o_x_15[1];
  assign uSystolicPE_254_io_clear_o = clear_o_x_15[1];
  assign ofm_x_15_0 = uSystolicPE_254_io_ofm_d;
  assign randW_x_0_16 = uSystolicPE_254_io_randW_d;
  assign uSystolicPEBorder_17_io_mac_done = mac_done_x_1[0];
  assign uSystolicPEBorder_17_io_enable_i = enable_i_x_1[0];
  assign uSystolicPEBorder_17_io_clear_i = clear_i_x_1[0];
  assign ifm_sign_x_1_1 = uSystolicPEBorder_17_io_ifm_sign_d;
  assign ifm_dff_x_1_1 = uSystolicPEBorder_17_io_ifm_dff_d;
  assign uSystolicPEBorder_17_io_enable_w = enable_w_x_0[1];
  assign uSystolicPEBorder_17_io_clear_w = clear_w_x_0[1];
  assign wght_sign_x_0_2 = uSystolicPEBorder_17_io_wght_sign_d;
  assign wght_abs_x_0_2 = uSystolicPEBorder_17_io_wght_abs_d;
  assign uSystolicPEBorder_17_io_enable_o = enable_o_x_0[2];
  assign uSystolicPEBorder_17_io_clear_o = clear_o_x_0[2];
  assign ofm_x_0_1 = uSystolicPEBorder_17_io_ofm_d;
  assign randW_x_1_1 = uSystolicPEBorder_17_io_randW_d;
  assign uSystolicPE_255_io_mac_done = mac_done_x_1[1];
  assign uSystolicPE_255_io_enable_i = enable_i_x_1[1];
  assign uSystolicPE_255_io_clear_i = clear_i_x_1[1];
  assign ifm_sign_x_1_2 = uSystolicPE_255_io_ifm_sign_d;
  assign ifm_dff_x_1_2 = uSystolicPE_255_io_ifm_dff_d;
  assign uSystolicPE_255_io_enable_w = enable_w_x_1[1];
  assign uSystolicPE_255_io_clear_w = clear_w_x_1[1];
  assign wght_sign_x_1_2 = uSystolicPE_255_io_wght_sign_d;
  assign wght_abs_x_1_2 = uSystolicPE_255_io_wght_abs_d;
  assign uSystolicPE_255_io_enable_o = enable_o_x_1[2];
  assign uSystolicPE_255_io_clear_o = clear_o_x_1[2];
  assign ofm_x_1_1 = uSystolicPE_255_io_ofm_d;
  assign randW_x_1_2 = uSystolicPE_255_io_randW_d;
  assign uSystolicPE_256_io_mac_done = mac_done_x_1[2];
  assign uSystolicPE_256_io_enable_i = enable_i_x_1[2];
  assign uSystolicPE_256_io_clear_i = clear_i_x_1[2];
  assign ifm_sign_x_1_3 = uSystolicPE_256_io_ifm_sign_d;
  assign ifm_dff_x_1_3 = uSystolicPE_256_io_ifm_dff_d;
  assign uSystolicPE_256_io_enable_w = enable_w_x_2[1];
  assign uSystolicPE_256_io_clear_w = clear_w_x_2[1];
  assign wght_sign_x_2_2 = uSystolicPE_256_io_wght_sign_d;
  assign wght_abs_x_2_2 = uSystolicPE_256_io_wght_abs_d;
  assign uSystolicPE_256_io_enable_o = enable_o_x_2[2];
  assign uSystolicPE_256_io_clear_o = clear_o_x_2[2];
  assign ofm_x_2_1 = uSystolicPE_256_io_ofm_d;
  assign randW_x_1_3 = uSystolicPE_256_io_randW_d;
  assign uSystolicPE_257_io_mac_done = mac_done_x_1[3];
  assign uSystolicPE_257_io_enable_i = enable_i_x_1[3];
  assign uSystolicPE_257_io_clear_i = clear_i_x_1[3];
  assign ifm_sign_x_1_4 = uSystolicPE_257_io_ifm_sign_d;
  assign ifm_dff_x_1_4 = uSystolicPE_257_io_ifm_dff_d;
  assign uSystolicPE_257_io_enable_w = enable_w_x_3[1];
  assign uSystolicPE_257_io_clear_w = clear_w_x_3[1];
  assign wght_sign_x_3_2 = uSystolicPE_257_io_wght_sign_d;
  assign wght_abs_x_3_2 = uSystolicPE_257_io_wght_abs_d;
  assign uSystolicPE_257_io_enable_o = enable_o_x_3[2];
  assign uSystolicPE_257_io_clear_o = clear_o_x_3[2];
  assign ofm_x_3_1 = uSystolicPE_257_io_ofm_d;
  assign randW_x_1_4 = uSystolicPE_257_io_randW_d;
  assign uSystolicPE_258_io_mac_done = mac_done_x_1[4];
  assign uSystolicPE_258_io_enable_i = enable_i_x_1[4];
  assign uSystolicPE_258_io_clear_i = clear_i_x_1[4];
  assign ifm_sign_x_1_5 = uSystolicPE_258_io_ifm_sign_d;
  assign ifm_dff_x_1_5 = uSystolicPE_258_io_ifm_dff_d;
  assign uSystolicPE_258_io_enable_w = enable_w_x_4[1];
  assign uSystolicPE_258_io_clear_w = clear_w_x_4[1];
  assign wght_sign_x_4_2 = uSystolicPE_258_io_wght_sign_d;
  assign wght_abs_x_4_2 = uSystolicPE_258_io_wght_abs_d;
  assign uSystolicPE_258_io_enable_o = enable_o_x_4[2];
  assign uSystolicPE_258_io_clear_o = clear_o_x_4[2];
  assign ofm_x_4_1 = uSystolicPE_258_io_ofm_d;
  assign randW_x_1_5 = uSystolicPE_258_io_randW_d;
  assign uSystolicPE_259_io_mac_done = mac_done_x_1[5];
  assign uSystolicPE_259_io_enable_i = enable_i_x_1[5];
  assign uSystolicPE_259_io_clear_i = clear_i_x_1[5];
  assign ifm_sign_x_1_6 = uSystolicPE_259_io_ifm_sign_d;
  assign ifm_dff_x_1_6 = uSystolicPE_259_io_ifm_dff_d;
  assign uSystolicPE_259_io_enable_w = enable_w_x_5[1];
  assign uSystolicPE_259_io_clear_w = clear_w_x_5[1];
  assign wght_sign_x_5_2 = uSystolicPE_259_io_wght_sign_d;
  assign wght_abs_x_5_2 = uSystolicPE_259_io_wght_abs_d;
  assign uSystolicPE_259_io_enable_o = enable_o_x_5[2];
  assign uSystolicPE_259_io_clear_o = clear_o_x_5[2];
  assign ofm_x_5_1 = uSystolicPE_259_io_ofm_d;
  assign randW_x_1_6 = uSystolicPE_259_io_randW_d;
  assign uSystolicPE_260_io_mac_done = mac_done_x_1[6];
  assign uSystolicPE_260_io_enable_i = enable_i_x_1[6];
  assign uSystolicPE_260_io_clear_i = clear_i_x_1[6];
  assign ifm_sign_x_1_7 = uSystolicPE_260_io_ifm_sign_d;
  assign ifm_dff_x_1_7 = uSystolicPE_260_io_ifm_dff_d;
  assign uSystolicPE_260_io_enable_w = enable_w_x_6[1];
  assign uSystolicPE_260_io_clear_w = clear_w_x_6[1];
  assign wght_sign_x_6_2 = uSystolicPE_260_io_wght_sign_d;
  assign wght_abs_x_6_2 = uSystolicPE_260_io_wght_abs_d;
  assign uSystolicPE_260_io_enable_o = enable_o_x_6[2];
  assign uSystolicPE_260_io_clear_o = clear_o_x_6[2];
  assign ofm_x_6_1 = uSystolicPE_260_io_ofm_d;
  assign randW_x_1_7 = uSystolicPE_260_io_randW_d;
  assign uSystolicPE_261_io_mac_done = mac_done_x_1[7];
  assign uSystolicPE_261_io_enable_i = enable_i_x_1[7];
  assign uSystolicPE_261_io_clear_i = clear_i_x_1[7];
  assign ifm_sign_x_1_8 = uSystolicPE_261_io_ifm_sign_d;
  assign ifm_dff_x_1_8 = uSystolicPE_261_io_ifm_dff_d;
  assign uSystolicPE_261_io_enable_w = enable_w_x_7[1];
  assign uSystolicPE_261_io_clear_w = clear_w_x_7[1];
  assign wght_sign_x_7_2 = uSystolicPE_261_io_wght_sign_d;
  assign wght_abs_x_7_2 = uSystolicPE_261_io_wght_abs_d;
  assign uSystolicPE_261_io_enable_o = enable_o_x_7[2];
  assign uSystolicPE_261_io_clear_o = clear_o_x_7[2];
  assign ofm_x_7_1 = uSystolicPE_261_io_ofm_d;
  assign randW_x_1_8 = uSystolicPE_261_io_randW_d;
  assign uSystolicPE_262_io_mac_done = mac_done_x_1[8];
  assign uSystolicPE_262_io_enable_i = enable_i_x_1[8];
  assign uSystolicPE_262_io_clear_i = clear_i_x_1[8];
  assign ifm_sign_x_1_9 = uSystolicPE_262_io_ifm_sign_d;
  assign ifm_dff_x_1_9 = uSystolicPE_262_io_ifm_dff_d;
  assign uSystolicPE_262_io_enable_w = enable_w_x_8[1];
  assign uSystolicPE_262_io_clear_w = clear_w_x_8[1];
  assign wght_sign_x_8_2 = uSystolicPE_262_io_wght_sign_d;
  assign wght_abs_x_8_2 = uSystolicPE_262_io_wght_abs_d;
  assign uSystolicPE_262_io_enable_o = enable_o_x_8[2];
  assign uSystolicPE_262_io_clear_o = clear_o_x_8[2];
  assign ofm_x_8_1 = uSystolicPE_262_io_ofm_d;
  assign randW_x_1_9 = uSystolicPE_262_io_randW_d;
  assign uSystolicPE_263_io_mac_done = mac_done_x_1[9];
  assign uSystolicPE_263_io_enable_i = enable_i_x_1[9];
  assign uSystolicPE_263_io_clear_i = clear_i_x_1[9];
  assign ifm_sign_x_1_10 = uSystolicPE_263_io_ifm_sign_d;
  assign ifm_dff_x_1_10 = uSystolicPE_263_io_ifm_dff_d;
  assign uSystolicPE_263_io_enable_w = enable_w_x_9[1];
  assign uSystolicPE_263_io_clear_w = clear_w_x_9[1];
  assign wght_sign_x_9_2 = uSystolicPE_263_io_wght_sign_d;
  assign wght_abs_x_9_2 = uSystolicPE_263_io_wght_abs_d;
  assign uSystolicPE_263_io_enable_o = enable_o_x_9[2];
  assign uSystolicPE_263_io_clear_o = clear_o_x_9[2];
  assign ofm_x_9_1 = uSystolicPE_263_io_ofm_d;
  assign randW_x_1_10 = uSystolicPE_263_io_randW_d;
  assign uSystolicPE_264_io_mac_done = mac_done_x_1[10];
  assign uSystolicPE_264_io_enable_i = enable_i_x_1[10];
  assign uSystolicPE_264_io_clear_i = clear_i_x_1[10];
  assign ifm_sign_x_1_11 = uSystolicPE_264_io_ifm_sign_d;
  assign ifm_dff_x_1_11 = uSystolicPE_264_io_ifm_dff_d;
  assign uSystolicPE_264_io_enable_w = enable_w_x_10[1];
  assign uSystolicPE_264_io_clear_w = clear_w_x_10[1];
  assign wght_sign_x_10_2 = uSystolicPE_264_io_wght_sign_d;
  assign wght_abs_x_10_2 = uSystolicPE_264_io_wght_abs_d;
  assign uSystolicPE_264_io_enable_o = enable_o_x_10[2];
  assign uSystolicPE_264_io_clear_o = clear_o_x_10[2];
  assign ofm_x_10_1 = uSystolicPE_264_io_ofm_d;
  assign randW_x_1_11 = uSystolicPE_264_io_randW_d;
  assign uSystolicPE_265_io_mac_done = mac_done_x_1[11];
  assign uSystolicPE_265_io_enable_i = enable_i_x_1[11];
  assign uSystolicPE_265_io_clear_i = clear_i_x_1[11];
  assign ifm_sign_x_1_12 = uSystolicPE_265_io_ifm_sign_d;
  assign ifm_dff_x_1_12 = uSystolicPE_265_io_ifm_dff_d;
  assign uSystolicPE_265_io_enable_w = enable_w_x_11[1];
  assign uSystolicPE_265_io_clear_w = clear_w_x_11[1];
  assign wght_sign_x_11_2 = uSystolicPE_265_io_wght_sign_d;
  assign wght_abs_x_11_2 = uSystolicPE_265_io_wght_abs_d;
  assign uSystolicPE_265_io_enable_o = enable_o_x_11[2];
  assign uSystolicPE_265_io_clear_o = clear_o_x_11[2];
  assign ofm_x_11_1 = uSystolicPE_265_io_ofm_d;
  assign randW_x_1_12 = uSystolicPE_265_io_randW_d;
  assign uSystolicPE_266_io_mac_done = mac_done_x_1[12];
  assign uSystolicPE_266_io_enable_i = enable_i_x_1[12];
  assign uSystolicPE_266_io_clear_i = clear_i_x_1[12];
  assign ifm_sign_x_1_13 = uSystolicPE_266_io_ifm_sign_d;
  assign ifm_dff_x_1_13 = uSystolicPE_266_io_ifm_dff_d;
  assign uSystolicPE_266_io_enable_w = enable_w_x_12[1];
  assign uSystolicPE_266_io_clear_w = clear_w_x_12[1];
  assign wght_sign_x_12_2 = uSystolicPE_266_io_wght_sign_d;
  assign wght_abs_x_12_2 = uSystolicPE_266_io_wght_abs_d;
  assign uSystolicPE_266_io_enable_o = enable_o_x_12[2];
  assign uSystolicPE_266_io_clear_o = clear_o_x_12[2];
  assign ofm_x_12_1 = uSystolicPE_266_io_ofm_d;
  assign randW_x_1_13 = uSystolicPE_266_io_randW_d;
  assign uSystolicPE_267_io_mac_done = mac_done_x_1[13];
  assign uSystolicPE_267_io_enable_i = enable_i_x_1[13];
  assign uSystolicPE_267_io_clear_i = clear_i_x_1[13];
  assign ifm_sign_x_1_14 = uSystolicPE_267_io_ifm_sign_d;
  assign ifm_dff_x_1_14 = uSystolicPE_267_io_ifm_dff_d;
  assign uSystolicPE_267_io_enable_w = enable_w_x_13[1];
  assign uSystolicPE_267_io_clear_w = clear_w_x_13[1];
  assign wght_sign_x_13_2 = uSystolicPE_267_io_wght_sign_d;
  assign wght_abs_x_13_2 = uSystolicPE_267_io_wght_abs_d;
  assign uSystolicPE_267_io_enable_o = enable_o_x_13[2];
  assign uSystolicPE_267_io_clear_o = clear_o_x_13[2];
  assign ofm_x_13_1 = uSystolicPE_267_io_ofm_d;
  assign randW_x_1_14 = uSystolicPE_267_io_randW_d;
  assign uSystolicPE_268_io_mac_done = mac_done_x_1[14];
  assign uSystolicPE_268_io_enable_i = enable_i_x_1[14];
  assign uSystolicPE_268_io_clear_i = clear_i_x_1[14];
  assign ifm_sign_x_1_15 = uSystolicPE_268_io_ifm_sign_d;
  assign ifm_dff_x_1_15 = uSystolicPE_268_io_ifm_dff_d;
  assign uSystolicPE_268_io_enable_w = enable_w_x_14[1];
  assign uSystolicPE_268_io_clear_w = clear_w_x_14[1];
  assign wght_sign_x_14_2 = uSystolicPE_268_io_wght_sign_d;
  assign wght_abs_x_14_2 = uSystolicPE_268_io_wght_abs_d;
  assign uSystolicPE_268_io_enable_o = enable_o_x_14[2];
  assign uSystolicPE_268_io_clear_o = clear_o_x_14[2];
  assign ofm_x_14_1 = uSystolicPE_268_io_ofm_d;
  assign randW_x_1_15 = uSystolicPE_268_io_randW_d;
  assign uSystolicPE_269_io_mac_done = mac_done_x_1[15];
  assign uSystolicPE_269_io_enable_i = enable_i_x_1[15];
  assign uSystolicPE_269_io_clear_i = clear_i_x_1[15];
  assign ifm_sign_x_1_16 = uSystolicPE_269_io_ifm_sign_d;
  assign ifm_dff_x_1_16 = uSystolicPE_269_io_ifm_dff_d;
  assign uSystolicPE_269_io_enable_w = enable_w_x_15[1];
  assign uSystolicPE_269_io_clear_w = clear_w_x_15[1];
  assign wght_sign_x_15_2 = uSystolicPE_269_io_wght_sign_d;
  assign wght_abs_x_15_2 = uSystolicPE_269_io_wght_abs_d;
  assign uSystolicPE_269_io_enable_o = enable_o_x_15[2];
  assign uSystolicPE_269_io_clear_o = clear_o_x_15[2];
  assign ofm_x_15_1 = uSystolicPE_269_io_ofm_d;
  assign randW_x_1_16 = uSystolicPE_269_io_randW_d;
  assign uSystolicPEBorder_18_io_mac_done = mac_done_x_2[0];
  assign uSystolicPEBorder_18_io_enable_i = enable_i_x_2[0];
  assign uSystolicPEBorder_18_io_clear_i = clear_i_x_2[0];
  assign ifm_sign_x_2_1 = uSystolicPEBorder_18_io_ifm_sign_d;
  assign ifm_dff_x_2_1 = uSystolicPEBorder_18_io_ifm_dff_d;
  assign uSystolicPEBorder_18_io_enable_w = enable_w_x_0[2];
  assign uSystolicPEBorder_18_io_clear_w = clear_w_x_0[2];
  assign wght_sign_x_0_3 = uSystolicPEBorder_18_io_wght_sign_d;
  assign wght_abs_x_0_3 = uSystolicPEBorder_18_io_wght_abs_d;
  assign uSystolicPEBorder_18_io_enable_o = enable_o_x_0[3];
  assign uSystolicPEBorder_18_io_clear_o = clear_o_x_0[3];
  assign ofm_x_0_2 = uSystolicPEBorder_18_io_ofm_d;
  assign randW_x_2_1 = uSystolicPEBorder_18_io_randW_d;
  assign uSystolicPE_270_io_mac_done = mac_done_x_2[1];
  assign uSystolicPE_270_io_enable_i = enable_i_x_2[1];
  assign uSystolicPE_270_io_clear_i = clear_i_x_2[1];
  assign ifm_sign_x_2_2 = uSystolicPE_270_io_ifm_sign_d;
  assign ifm_dff_x_2_2 = uSystolicPE_270_io_ifm_dff_d;
  assign uSystolicPE_270_io_enable_w = enable_w_x_1[2];
  assign uSystolicPE_270_io_clear_w = clear_w_x_1[2];
  assign wght_sign_x_1_3 = uSystolicPE_270_io_wght_sign_d;
  assign wght_abs_x_1_3 = uSystolicPE_270_io_wght_abs_d;
  assign uSystolicPE_270_io_enable_o = enable_o_x_1[3];
  assign uSystolicPE_270_io_clear_o = clear_o_x_1[3];
  assign ofm_x_1_2 = uSystolicPE_270_io_ofm_d;
  assign randW_x_2_2 = uSystolicPE_270_io_randW_d;
  assign uSystolicPE_271_io_mac_done = mac_done_x_2[2];
  assign uSystolicPE_271_io_enable_i = enable_i_x_2[2];
  assign uSystolicPE_271_io_clear_i = clear_i_x_2[2];
  assign ifm_sign_x_2_3 = uSystolicPE_271_io_ifm_sign_d;
  assign ifm_dff_x_2_3 = uSystolicPE_271_io_ifm_dff_d;
  assign uSystolicPE_271_io_enable_w = enable_w_x_2[2];
  assign uSystolicPE_271_io_clear_w = clear_w_x_2[2];
  assign wght_sign_x_2_3 = uSystolicPE_271_io_wght_sign_d;
  assign wght_abs_x_2_3 = uSystolicPE_271_io_wght_abs_d;
  assign uSystolicPE_271_io_enable_o = enable_o_x_2[3];
  assign uSystolicPE_271_io_clear_o = clear_o_x_2[3];
  assign ofm_x_2_2 = uSystolicPE_271_io_ofm_d;
  assign randW_x_2_3 = uSystolicPE_271_io_randW_d;
  assign uSystolicPE_272_io_mac_done = mac_done_x_2[3];
  assign uSystolicPE_272_io_enable_i = enable_i_x_2[3];
  assign uSystolicPE_272_io_clear_i = clear_i_x_2[3];
  assign ifm_sign_x_2_4 = uSystolicPE_272_io_ifm_sign_d;
  assign ifm_dff_x_2_4 = uSystolicPE_272_io_ifm_dff_d;
  assign uSystolicPE_272_io_enable_w = enable_w_x_3[2];
  assign uSystolicPE_272_io_clear_w = clear_w_x_3[2];
  assign wght_sign_x_3_3 = uSystolicPE_272_io_wght_sign_d;
  assign wght_abs_x_3_3 = uSystolicPE_272_io_wght_abs_d;
  assign uSystolicPE_272_io_enable_o = enable_o_x_3[3];
  assign uSystolicPE_272_io_clear_o = clear_o_x_3[3];
  assign ofm_x_3_2 = uSystolicPE_272_io_ofm_d;
  assign randW_x_2_4 = uSystolicPE_272_io_randW_d;
  assign uSystolicPE_273_io_mac_done = mac_done_x_2[4];
  assign uSystolicPE_273_io_enable_i = enable_i_x_2[4];
  assign uSystolicPE_273_io_clear_i = clear_i_x_2[4];
  assign ifm_sign_x_2_5 = uSystolicPE_273_io_ifm_sign_d;
  assign ifm_dff_x_2_5 = uSystolicPE_273_io_ifm_dff_d;
  assign uSystolicPE_273_io_enable_w = enable_w_x_4[2];
  assign uSystolicPE_273_io_clear_w = clear_w_x_4[2];
  assign wght_sign_x_4_3 = uSystolicPE_273_io_wght_sign_d;
  assign wght_abs_x_4_3 = uSystolicPE_273_io_wght_abs_d;
  assign uSystolicPE_273_io_enable_o = enable_o_x_4[3];
  assign uSystolicPE_273_io_clear_o = clear_o_x_4[3];
  assign ofm_x_4_2 = uSystolicPE_273_io_ofm_d;
  assign randW_x_2_5 = uSystolicPE_273_io_randW_d;
  assign uSystolicPE_274_io_mac_done = mac_done_x_2[5];
  assign uSystolicPE_274_io_enable_i = enable_i_x_2[5];
  assign uSystolicPE_274_io_clear_i = clear_i_x_2[5];
  assign ifm_sign_x_2_6 = uSystolicPE_274_io_ifm_sign_d;
  assign ifm_dff_x_2_6 = uSystolicPE_274_io_ifm_dff_d;
  assign uSystolicPE_274_io_enable_w = enable_w_x_5[2];
  assign uSystolicPE_274_io_clear_w = clear_w_x_5[2];
  assign wght_sign_x_5_3 = uSystolicPE_274_io_wght_sign_d;
  assign wght_abs_x_5_3 = uSystolicPE_274_io_wght_abs_d;
  assign uSystolicPE_274_io_enable_o = enable_o_x_5[3];
  assign uSystolicPE_274_io_clear_o = clear_o_x_5[3];
  assign ofm_x_5_2 = uSystolicPE_274_io_ofm_d;
  assign randW_x_2_6 = uSystolicPE_274_io_randW_d;
  assign uSystolicPE_275_io_mac_done = mac_done_x_2[6];
  assign uSystolicPE_275_io_enable_i = enable_i_x_2[6];
  assign uSystolicPE_275_io_clear_i = clear_i_x_2[6];
  assign ifm_sign_x_2_7 = uSystolicPE_275_io_ifm_sign_d;
  assign ifm_dff_x_2_7 = uSystolicPE_275_io_ifm_dff_d;
  assign uSystolicPE_275_io_enable_w = enable_w_x_6[2];
  assign uSystolicPE_275_io_clear_w = clear_w_x_6[2];
  assign wght_sign_x_6_3 = uSystolicPE_275_io_wght_sign_d;
  assign wght_abs_x_6_3 = uSystolicPE_275_io_wght_abs_d;
  assign uSystolicPE_275_io_enable_o = enable_o_x_6[3];
  assign uSystolicPE_275_io_clear_o = clear_o_x_6[3];
  assign ofm_x_6_2 = uSystolicPE_275_io_ofm_d;
  assign randW_x_2_7 = uSystolicPE_275_io_randW_d;
  assign uSystolicPE_276_io_mac_done = mac_done_x_2[7];
  assign uSystolicPE_276_io_enable_i = enable_i_x_2[7];
  assign uSystolicPE_276_io_clear_i = clear_i_x_2[7];
  assign ifm_sign_x_2_8 = uSystolicPE_276_io_ifm_sign_d;
  assign ifm_dff_x_2_8 = uSystolicPE_276_io_ifm_dff_d;
  assign uSystolicPE_276_io_enable_w = enable_w_x_7[2];
  assign uSystolicPE_276_io_clear_w = clear_w_x_7[2];
  assign wght_sign_x_7_3 = uSystolicPE_276_io_wght_sign_d;
  assign wght_abs_x_7_3 = uSystolicPE_276_io_wght_abs_d;
  assign uSystolicPE_276_io_enable_o = enable_o_x_7[3];
  assign uSystolicPE_276_io_clear_o = clear_o_x_7[3];
  assign ofm_x_7_2 = uSystolicPE_276_io_ofm_d;
  assign randW_x_2_8 = uSystolicPE_276_io_randW_d;
  assign uSystolicPE_277_io_mac_done = mac_done_x_2[8];
  assign uSystolicPE_277_io_enable_i = enable_i_x_2[8];
  assign uSystolicPE_277_io_clear_i = clear_i_x_2[8];
  assign ifm_sign_x_2_9 = uSystolicPE_277_io_ifm_sign_d;
  assign ifm_dff_x_2_9 = uSystolicPE_277_io_ifm_dff_d;
  assign uSystolicPE_277_io_enable_w = enable_w_x_8[2];
  assign uSystolicPE_277_io_clear_w = clear_w_x_8[2];
  assign wght_sign_x_8_3 = uSystolicPE_277_io_wght_sign_d;
  assign wght_abs_x_8_3 = uSystolicPE_277_io_wght_abs_d;
  assign uSystolicPE_277_io_enable_o = enable_o_x_8[3];
  assign uSystolicPE_277_io_clear_o = clear_o_x_8[3];
  assign ofm_x_8_2 = uSystolicPE_277_io_ofm_d;
  assign randW_x_2_9 = uSystolicPE_277_io_randW_d;
  assign uSystolicPE_278_io_mac_done = mac_done_x_2[9];
  assign uSystolicPE_278_io_enable_i = enable_i_x_2[9];
  assign uSystolicPE_278_io_clear_i = clear_i_x_2[9];
  assign ifm_sign_x_2_10 = uSystolicPE_278_io_ifm_sign_d;
  assign ifm_dff_x_2_10 = uSystolicPE_278_io_ifm_dff_d;
  assign uSystolicPE_278_io_enable_w = enable_w_x_9[2];
  assign uSystolicPE_278_io_clear_w = clear_w_x_9[2];
  assign wght_sign_x_9_3 = uSystolicPE_278_io_wght_sign_d;
  assign wght_abs_x_9_3 = uSystolicPE_278_io_wght_abs_d;
  assign uSystolicPE_278_io_enable_o = enable_o_x_9[3];
  assign uSystolicPE_278_io_clear_o = clear_o_x_9[3];
  assign ofm_x_9_2 = uSystolicPE_278_io_ofm_d;
  assign randW_x_2_10 = uSystolicPE_278_io_randW_d;
  assign uSystolicPE_279_io_mac_done = mac_done_x_2[10];
  assign uSystolicPE_279_io_enable_i = enable_i_x_2[10];
  assign uSystolicPE_279_io_clear_i = clear_i_x_2[10];
  assign ifm_sign_x_2_11 = uSystolicPE_279_io_ifm_sign_d;
  assign ifm_dff_x_2_11 = uSystolicPE_279_io_ifm_dff_d;
  assign uSystolicPE_279_io_enable_w = enable_w_x_10[2];
  assign uSystolicPE_279_io_clear_w = clear_w_x_10[2];
  assign wght_sign_x_10_3 = uSystolicPE_279_io_wght_sign_d;
  assign wght_abs_x_10_3 = uSystolicPE_279_io_wght_abs_d;
  assign uSystolicPE_279_io_enable_o = enable_o_x_10[3];
  assign uSystolicPE_279_io_clear_o = clear_o_x_10[3];
  assign ofm_x_10_2 = uSystolicPE_279_io_ofm_d;
  assign randW_x_2_11 = uSystolicPE_279_io_randW_d;
  assign uSystolicPE_280_io_mac_done = mac_done_x_2[11];
  assign uSystolicPE_280_io_enable_i = enable_i_x_2[11];
  assign uSystolicPE_280_io_clear_i = clear_i_x_2[11];
  assign ifm_sign_x_2_12 = uSystolicPE_280_io_ifm_sign_d;
  assign ifm_dff_x_2_12 = uSystolicPE_280_io_ifm_dff_d;
  assign uSystolicPE_280_io_enable_w = enable_w_x_11[2];
  assign uSystolicPE_280_io_clear_w = clear_w_x_11[2];
  assign wght_sign_x_11_3 = uSystolicPE_280_io_wght_sign_d;
  assign wght_abs_x_11_3 = uSystolicPE_280_io_wght_abs_d;
  assign uSystolicPE_280_io_enable_o = enable_o_x_11[3];
  assign uSystolicPE_280_io_clear_o = clear_o_x_11[3];
  assign ofm_x_11_2 = uSystolicPE_280_io_ofm_d;
  assign randW_x_2_12 = uSystolicPE_280_io_randW_d;
  assign uSystolicPE_281_io_mac_done = mac_done_x_2[12];
  assign uSystolicPE_281_io_enable_i = enable_i_x_2[12];
  assign uSystolicPE_281_io_clear_i = clear_i_x_2[12];
  assign ifm_sign_x_2_13 = uSystolicPE_281_io_ifm_sign_d;
  assign ifm_dff_x_2_13 = uSystolicPE_281_io_ifm_dff_d;
  assign uSystolicPE_281_io_enable_w = enable_w_x_12[2];
  assign uSystolicPE_281_io_clear_w = clear_w_x_12[2];
  assign wght_sign_x_12_3 = uSystolicPE_281_io_wght_sign_d;
  assign wght_abs_x_12_3 = uSystolicPE_281_io_wght_abs_d;
  assign uSystolicPE_281_io_enable_o = enable_o_x_12[3];
  assign uSystolicPE_281_io_clear_o = clear_o_x_12[3];
  assign ofm_x_12_2 = uSystolicPE_281_io_ofm_d;
  assign randW_x_2_13 = uSystolicPE_281_io_randW_d;
  assign uSystolicPE_282_io_mac_done = mac_done_x_2[13];
  assign uSystolicPE_282_io_enable_i = enable_i_x_2[13];
  assign uSystolicPE_282_io_clear_i = clear_i_x_2[13];
  assign ifm_sign_x_2_14 = uSystolicPE_282_io_ifm_sign_d;
  assign ifm_dff_x_2_14 = uSystolicPE_282_io_ifm_dff_d;
  assign uSystolicPE_282_io_enable_w = enable_w_x_13[2];
  assign uSystolicPE_282_io_clear_w = clear_w_x_13[2];
  assign wght_sign_x_13_3 = uSystolicPE_282_io_wght_sign_d;
  assign wght_abs_x_13_3 = uSystolicPE_282_io_wght_abs_d;
  assign uSystolicPE_282_io_enable_o = enable_o_x_13[3];
  assign uSystolicPE_282_io_clear_o = clear_o_x_13[3];
  assign ofm_x_13_2 = uSystolicPE_282_io_ofm_d;
  assign randW_x_2_14 = uSystolicPE_282_io_randW_d;
  assign uSystolicPE_283_io_mac_done = mac_done_x_2[14];
  assign uSystolicPE_283_io_enable_i = enable_i_x_2[14];
  assign uSystolicPE_283_io_clear_i = clear_i_x_2[14];
  assign ifm_sign_x_2_15 = uSystolicPE_283_io_ifm_sign_d;
  assign ifm_dff_x_2_15 = uSystolicPE_283_io_ifm_dff_d;
  assign uSystolicPE_283_io_enable_w = enable_w_x_14[2];
  assign uSystolicPE_283_io_clear_w = clear_w_x_14[2];
  assign wght_sign_x_14_3 = uSystolicPE_283_io_wght_sign_d;
  assign wght_abs_x_14_3 = uSystolicPE_283_io_wght_abs_d;
  assign uSystolicPE_283_io_enable_o = enable_o_x_14[3];
  assign uSystolicPE_283_io_clear_o = clear_o_x_14[3];
  assign ofm_x_14_2 = uSystolicPE_283_io_ofm_d;
  assign randW_x_2_15 = uSystolicPE_283_io_randW_d;
  assign uSystolicPE_284_io_mac_done = mac_done_x_2[15];
  assign uSystolicPE_284_io_enable_i = enable_i_x_2[15];
  assign uSystolicPE_284_io_clear_i = clear_i_x_2[15];
  assign ifm_sign_x_2_16 = uSystolicPE_284_io_ifm_sign_d;
  assign ifm_dff_x_2_16 = uSystolicPE_284_io_ifm_dff_d;
  assign uSystolicPE_284_io_enable_w = enable_w_x_15[2];
  assign uSystolicPE_284_io_clear_w = clear_w_x_15[2];
  assign wght_sign_x_15_3 = uSystolicPE_284_io_wght_sign_d;
  assign wght_abs_x_15_3 = uSystolicPE_284_io_wght_abs_d;
  assign uSystolicPE_284_io_enable_o = enable_o_x_15[3];
  assign uSystolicPE_284_io_clear_o = clear_o_x_15[3];
  assign ofm_x_15_2 = uSystolicPE_284_io_ofm_d;
  assign randW_x_2_16 = uSystolicPE_284_io_randW_d;
  assign uSystolicPEBorder_19_io_mac_done = mac_done_x_3[0];
  assign uSystolicPEBorder_19_io_enable_i = enable_i_x_3[0];
  assign uSystolicPEBorder_19_io_clear_i = clear_i_x_3[0];
  assign ifm_sign_x_3_1 = uSystolicPEBorder_19_io_ifm_sign_d;
  assign ifm_dff_x_3_1 = uSystolicPEBorder_19_io_ifm_dff_d;
  assign uSystolicPEBorder_19_io_enable_w = enable_w_x_0[3];
  assign uSystolicPEBorder_19_io_clear_w = clear_w_x_0[3];
  assign wght_sign_x_0_4 = uSystolicPEBorder_19_io_wght_sign_d;
  assign wght_abs_x_0_4 = uSystolicPEBorder_19_io_wght_abs_d;
  assign uSystolicPEBorder_19_io_enable_o = enable_o_x_0[4];
  assign uSystolicPEBorder_19_io_clear_o = clear_o_x_0[4];
  assign ofm_x_0_3 = uSystolicPEBorder_19_io_ofm_d;
  assign randW_x_3_1 = uSystolicPEBorder_19_io_randW_d;
  assign uSystolicPE_285_io_mac_done = mac_done_x_3[1];
  assign uSystolicPE_285_io_enable_i = enable_i_x_3[1];
  assign uSystolicPE_285_io_clear_i = clear_i_x_3[1];
  assign ifm_sign_x_3_2 = uSystolicPE_285_io_ifm_sign_d;
  assign ifm_dff_x_3_2 = uSystolicPE_285_io_ifm_dff_d;
  assign uSystolicPE_285_io_enable_w = enable_w_x_1[3];
  assign uSystolicPE_285_io_clear_w = clear_w_x_1[3];
  assign wght_sign_x_1_4 = uSystolicPE_285_io_wght_sign_d;
  assign wght_abs_x_1_4 = uSystolicPE_285_io_wght_abs_d;
  assign uSystolicPE_285_io_enable_o = enable_o_x_1[4];
  assign uSystolicPE_285_io_clear_o = clear_o_x_1[4];
  assign ofm_x_1_3 = uSystolicPE_285_io_ofm_d;
  assign randW_x_3_2 = uSystolicPE_285_io_randW_d;
  assign uSystolicPE_286_io_mac_done = mac_done_x_3[2];
  assign uSystolicPE_286_io_enable_i = enable_i_x_3[2];
  assign uSystolicPE_286_io_clear_i = clear_i_x_3[2];
  assign ifm_sign_x_3_3 = uSystolicPE_286_io_ifm_sign_d;
  assign ifm_dff_x_3_3 = uSystolicPE_286_io_ifm_dff_d;
  assign uSystolicPE_286_io_enable_w = enable_w_x_2[3];
  assign uSystolicPE_286_io_clear_w = clear_w_x_2[3];
  assign wght_sign_x_2_4 = uSystolicPE_286_io_wght_sign_d;
  assign wght_abs_x_2_4 = uSystolicPE_286_io_wght_abs_d;
  assign uSystolicPE_286_io_enable_o = enable_o_x_2[4];
  assign uSystolicPE_286_io_clear_o = clear_o_x_2[4];
  assign ofm_x_2_3 = uSystolicPE_286_io_ofm_d;
  assign randW_x_3_3 = uSystolicPE_286_io_randW_d;
  assign uSystolicPE_287_io_mac_done = mac_done_x_3[3];
  assign uSystolicPE_287_io_enable_i = enable_i_x_3[3];
  assign uSystolicPE_287_io_clear_i = clear_i_x_3[3];
  assign ifm_sign_x_3_4 = uSystolicPE_287_io_ifm_sign_d;
  assign ifm_dff_x_3_4 = uSystolicPE_287_io_ifm_dff_d;
  assign uSystolicPE_287_io_enable_w = enable_w_x_3[3];
  assign uSystolicPE_287_io_clear_w = clear_w_x_3[3];
  assign wght_sign_x_3_4 = uSystolicPE_287_io_wght_sign_d;
  assign wght_abs_x_3_4 = uSystolicPE_287_io_wght_abs_d;
  assign uSystolicPE_287_io_enable_o = enable_o_x_3[4];
  assign uSystolicPE_287_io_clear_o = clear_o_x_3[4];
  assign ofm_x_3_3 = uSystolicPE_287_io_ofm_d;
  assign randW_x_3_4 = uSystolicPE_287_io_randW_d;
  assign uSystolicPE_288_io_mac_done = mac_done_x_3[4];
  assign uSystolicPE_288_io_enable_i = enable_i_x_3[4];
  assign uSystolicPE_288_io_clear_i = clear_i_x_3[4];
  assign ifm_sign_x_3_5 = uSystolicPE_288_io_ifm_sign_d;
  assign ifm_dff_x_3_5 = uSystolicPE_288_io_ifm_dff_d;
  assign uSystolicPE_288_io_enable_w = enable_w_x_4[3];
  assign uSystolicPE_288_io_clear_w = clear_w_x_4[3];
  assign wght_sign_x_4_4 = uSystolicPE_288_io_wght_sign_d;
  assign wght_abs_x_4_4 = uSystolicPE_288_io_wght_abs_d;
  assign uSystolicPE_288_io_enable_o = enable_o_x_4[4];
  assign uSystolicPE_288_io_clear_o = clear_o_x_4[4];
  assign ofm_x_4_3 = uSystolicPE_288_io_ofm_d;
  assign randW_x_3_5 = uSystolicPE_288_io_randW_d;
  assign uSystolicPE_289_io_mac_done = mac_done_x_3[5];
  assign uSystolicPE_289_io_enable_i = enable_i_x_3[5];
  assign uSystolicPE_289_io_clear_i = clear_i_x_3[5];
  assign ifm_sign_x_3_6 = uSystolicPE_289_io_ifm_sign_d;
  assign ifm_dff_x_3_6 = uSystolicPE_289_io_ifm_dff_d;
  assign uSystolicPE_289_io_enable_w = enable_w_x_5[3];
  assign uSystolicPE_289_io_clear_w = clear_w_x_5[3];
  assign wght_sign_x_5_4 = uSystolicPE_289_io_wght_sign_d;
  assign wght_abs_x_5_4 = uSystolicPE_289_io_wght_abs_d;
  assign uSystolicPE_289_io_enable_o = enable_o_x_5[4];
  assign uSystolicPE_289_io_clear_o = clear_o_x_5[4];
  assign ofm_x_5_3 = uSystolicPE_289_io_ofm_d;
  assign randW_x_3_6 = uSystolicPE_289_io_randW_d;
  assign uSystolicPE_290_io_mac_done = mac_done_x_3[6];
  assign uSystolicPE_290_io_enable_i = enable_i_x_3[6];
  assign uSystolicPE_290_io_clear_i = clear_i_x_3[6];
  assign ifm_sign_x_3_7 = uSystolicPE_290_io_ifm_sign_d;
  assign ifm_dff_x_3_7 = uSystolicPE_290_io_ifm_dff_d;
  assign uSystolicPE_290_io_enable_w = enable_w_x_6[3];
  assign uSystolicPE_290_io_clear_w = clear_w_x_6[3];
  assign wght_sign_x_6_4 = uSystolicPE_290_io_wght_sign_d;
  assign wght_abs_x_6_4 = uSystolicPE_290_io_wght_abs_d;
  assign uSystolicPE_290_io_enable_o = enable_o_x_6[4];
  assign uSystolicPE_290_io_clear_o = clear_o_x_6[4];
  assign ofm_x_6_3 = uSystolicPE_290_io_ofm_d;
  assign randW_x_3_7 = uSystolicPE_290_io_randW_d;
  assign uSystolicPE_291_io_mac_done = mac_done_x_3[7];
  assign uSystolicPE_291_io_enable_i = enable_i_x_3[7];
  assign uSystolicPE_291_io_clear_i = clear_i_x_3[7];
  assign ifm_sign_x_3_8 = uSystolicPE_291_io_ifm_sign_d;
  assign ifm_dff_x_3_8 = uSystolicPE_291_io_ifm_dff_d;
  assign uSystolicPE_291_io_enable_w = enable_w_x_7[3];
  assign uSystolicPE_291_io_clear_w = clear_w_x_7[3];
  assign wght_sign_x_7_4 = uSystolicPE_291_io_wght_sign_d;
  assign wght_abs_x_7_4 = uSystolicPE_291_io_wght_abs_d;
  assign uSystolicPE_291_io_enable_o = enable_o_x_7[4];
  assign uSystolicPE_291_io_clear_o = clear_o_x_7[4];
  assign ofm_x_7_3 = uSystolicPE_291_io_ofm_d;
  assign randW_x_3_8 = uSystolicPE_291_io_randW_d;
  assign uSystolicPE_292_io_mac_done = mac_done_x_3[8];
  assign uSystolicPE_292_io_enable_i = enable_i_x_3[8];
  assign uSystolicPE_292_io_clear_i = clear_i_x_3[8];
  assign ifm_sign_x_3_9 = uSystolicPE_292_io_ifm_sign_d;
  assign ifm_dff_x_3_9 = uSystolicPE_292_io_ifm_dff_d;
  assign uSystolicPE_292_io_enable_w = enable_w_x_8[3];
  assign uSystolicPE_292_io_clear_w = clear_w_x_8[3];
  assign wght_sign_x_8_4 = uSystolicPE_292_io_wght_sign_d;
  assign wght_abs_x_8_4 = uSystolicPE_292_io_wght_abs_d;
  assign uSystolicPE_292_io_enable_o = enable_o_x_8[4];
  assign uSystolicPE_292_io_clear_o = clear_o_x_8[4];
  assign ofm_x_8_3 = uSystolicPE_292_io_ofm_d;
  assign randW_x_3_9 = uSystolicPE_292_io_randW_d;
  assign uSystolicPE_293_io_mac_done = mac_done_x_3[9];
  assign uSystolicPE_293_io_enable_i = enable_i_x_3[9];
  assign uSystolicPE_293_io_clear_i = clear_i_x_3[9];
  assign ifm_sign_x_3_10 = uSystolicPE_293_io_ifm_sign_d;
  assign ifm_dff_x_3_10 = uSystolicPE_293_io_ifm_dff_d;
  assign uSystolicPE_293_io_enable_w = enable_w_x_9[3];
  assign uSystolicPE_293_io_clear_w = clear_w_x_9[3];
  assign wght_sign_x_9_4 = uSystolicPE_293_io_wght_sign_d;
  assign wght_abs_x_9_4 = uSystolicPE_293_io_wght_abs_d;
  assign uSystolicPE_293_io_enable_o = enable_o_x_9[4];
  assign uSystolicPE_293_io_clear_o = clear_o_x_9[4];
  assign ofm_x_9_3 = uSystolicPE_293_io_ofm_d;
  assign randW_x_3_10 = uSystolicPE_293_io_randW_d;
  assign uSystolicPE_294_io_mac_done = mac_done_x_3[10];
  assign uSystolicPE_294_io_enable_i = enable_i_x_3[10];
  assign uSystolicPE_294_io_clear_i = clear_i_x_3[10];
  assign ifm_sign_x_3_11 = uSystolicPE_294_io_ifm_sign_d;
  assign ifm_dff_x_3_11 = uSystolicPE_294_io_ifm_dff_d;
  assign uSystolicPE_294_io_enable_w = enable_w_x_10[3];
  assign uSystolicPE_294_io_clear_w = clear_w_x_10[3];
  assign wght_sign_x_10_4 = uSystolicPE_294_io_wght_sign_d;
  assign wght_abs_x_10_4 = uSystolicPE_294_io_wght_abs_d;
  assign uSystolicPE_294_io_enable_o = enable_o_x_10[4];
  assign uSystolicPE_294_io_clear_o = clear_o_x_10[4];
  assign ofm_x_10_3 = uSystolicPE_294_io_ofm_d;
  assign randW_x_3_11 = uSystolicPE_294_io_randW_d;
  assign uSystolicPE_295_io_mac_done = mac_done_x_3[11];
  assign uSystolicPE_295_io_enable_i = enable_i_x_3[11];
  assign uSystolicPE_295_io_clear_i = clear_i_x_3[11];
  assign ifm_sign_x_3_12 = uSystolicPE_295_io_ifm_sign_d;
  assign ifm_dff_x_3_12 = uSystolicPE_295_io_ifm_dff_d;
  assign uSystolicPE_295_io_enable_w = enable_w_x_11[3];
  assign uSystolicPE_295_io_clear_w = clear_w_x_11[3];
  assign wght_sign_x_11_4 = uSystolicPE_295_io_wght_sign_d;
  assign wght_abs_x_11_4 = uSystolicPE_295_io_wght_abs_d;
  assign uSystolicPE_295_io_enable_o = enable_o_x_11[4];
  assign uSystolicPE_295_io_clear_o = clear_o_x_11[4];
  assign ofm_x_11_3 = uSystolicPE_295_io_ofm_d;
  assign randW_x_3_12 = uSystolicPE_295_io_randW_d;
  assign uSystolicPE_296_io_mac_done = mac_done_x_3[12];
  assign uSystolicPE_296_io_enable_i = enable_i_x_3[12];
  assign uSystolicPE_296_io_clear_i = clear_i_x_3[12];
  assign ifm_sign_x_3_13 = uSystolicPE_296_io_ifm_sign_d;
  assign ifm_dff_x_3_13 = uSystolicPE_296_io_ifm_dff_d;
  assign uSystolicPE_296_io_enable_w = enable_w_x_12[3];
  assign uSystolicPE_296_io_clear_w = clear_w_x_12[3];
  assign wght_sign_x_12_4 = uSystolicPE_296_io_wght_sign_d;
  assign wght_abs_x_12_4 = uSystolicPE_296_io_wght_abs_d;
  assign uSystolicPE_296_io_enable_o = enable_o_x_12[4];
  assign uSystolicPE_296_io_clear_o = clear_o_x_12[4];
  assign ofm_x_12_3 = uSystolicPE_296_io_ofm_d;
  assign randW_x_3_13 = uSystolicPE_296_io_randW_d;
  assign uSystolicPE_297_io_mac_done = mac_done_x_3[13];
  assign uSystolicPE_297_io_enable_i = enable_i_x_3[13];
  assign uSystolicPE_297_io_clear_i = clear_i_x_3[13];
  assign ifm_sign_x_3_14 = uSystolicPE_297_io_ifm_sign_d;
  assign ifm_dff_x_3_14 = uSystolicPE_297_io_ifm_dff_d;
  assign uSystolicPE_297_io_enable_w = enable_w_x_13[3];
  assign uSystolicPE_297_io_clear_w = clear_w_x_13[3];
  assign wght_sign_x_13_4 = uSystolicPE_297_io_wght_sign_d;
  assign wght_abs_x_13_4 = uSystolicPE_297_io_wght_abs_d;
  assign uSystolicPE_297_io_enable_o = enable_o_x_13[4];
  assign uSystolicPE_297_io_clear_o = clear_o_x_13[4];
  assign ofm_x_13_3 = uSystolicPE_297_io_ofm_d;
  assign randW_x_3_14 = uSystolicPE_297_io_randW_d;
  assign uSystolicPE_298_io_mac_done = mac_done_x_3[14];
  assign uSystolicPE_298_io_enable_i = enable_i_x_3[14];
  assign uSystolicPE_298_io_clear_i = clear_i_x_3[14];
  assign ifm_sign_x_3_15 = uSystolicPE_298_io_ifm_sign_d;
  assign ifm_dff_x_3_15 = uSystolicPE_298_io_ifm_dff_d;
  assign uSystolicPE_298_io_enable_w = enable_w_x_14[3];
  assign uSystolicPE_298_io_clear_w = clear_w_x_14[3];
  assign wght_sign_x_14_4 = uSystolicPE_298_io_wght_sign_d;
  assign wght_abs_x_14_4 = uSystolicPE_298_io_wght_abs_d;
  assign uSystolicPE_298_io_enable_o = enable_o_x_14[4];
  assign uSystolicPE_298_io_clear_o = clear_o_x_14[4];
  assign ofm_x_14_3 = uSystolicPE_298_io_ofm_d;
  assign randW_x_3_15 = uSystolicPE_298_io_randW_d;
  assign uSystolicPE_299_io_mac_done = mac_done_x_3[15];
  assign uSystolicPE_299_io_enable_i = enable_i_x_3[15];
  assign uSystolicPE_299_io_clear_i = clear_i_x_3[15];
  assign ifm_sign_x_3_16 = uSystolicPE_299_io_ifm_sign_d;
  assign ifm_dff_x_3_16 = uSystolicPE_299_io_ifm_dff_d;
  assign uSystolicPE_299_io_enable_w = enable_w_x_15[3];
  assign uSystolicPE_299_io_clear_w = clear_w_x_15[3];
  assign wght_sign_x_15_4 = uSystolicPE_299_io_wght_sign_d;
  assign wght_abs_x_15_4 = uSystolicPE_299_io_wght_abs_d;
  assign uSystolicPE_299_io_enable_o = enable_o_x_15[4];
  assign uSystolicPE_299_io_clear_o = clear_o_x_15[4];
  assign ofm_x_15_3 = uSystolicPE_299_io_ofm_d;
  assign randW_x_3_16 = uSystolicPE_299_io_randW_d;
  assign uSystolicPEBorder_20_io_mac_done = mac_done_x_4[0];
  assign uSystolicPEBorder_20_io_enable_i = enable_i_x_4[0];
  assign uSystolicPEBorder_20_io_clear_i = clear_i_x_4[0];
  assign ifm_sign_x_4_1 = uSystolicPEBorder_20_io_ifm_sign_d;
  assign ifm_dff_x_4_1 = uSystolicPEBorder_20_io_ifm_dff_d;
  assign uSystolicPEBorder_20_io_enable_w = enable_w_x_0[4];
  assign uSystolicPEBorder_20_io_clear_w = clear_w_x_0[4];
  assign wght_sign_x_0_5 = uSystolicPEBorder_20_io_wght_sign_d;
  assign wght_abs_x_0_5 = uSystolicPEBorder_20_io_wght_abs_d;
  assign uSystolicPEBorder_20_io_enable_o = enable_o_x_0[5];
  assign uSystolicPEBorder_20_io_clear_o = clear_o_x_0[5];
  assign ofm_x_0_4 = uSystolicPEBorder_20_io_ofm_d;
  assign randW_x_4_1 = uSystolicPEBorder_20_io_randW_d;
  assign uSystolicPE_300_io_mac_done = mac_done_x_4[1];
  assign uSystolicPE_300_io_enable_i = enable_i_x_4[1];
  assign uSystolicPE_300_io_clear_i = clear_i_x_4[1];
  assign ifm_sign_x_4_2 = uSystolicPE_300_io_ifm_sign_d;
  assign ifm_dff_x_4_2 = uSystolicPE_300_io_ifm_dff_d;
  assign uSystolicPE_300_io_enable_w = enable_w_x_1[4];
  assign uSystolicPE_300_io_clear_w = clear_w_x_1[4];
  assign wght_sign_x_1_5 = uSystolicPE_300_io_wght_sign_d;
  assign wght_abs_x_1_5 = uSystolicPE_300_io_wght_abs_d;
  assign uSystolicPE_300_io_enable_o = enable_o_x_1[5];
  assign uSystolicPE_300_io_clear_o = clear_o_x_1[5];
  assign ofm_x_1_4 = uSystolicPE_300_io_ofm_d;
  assign randW_x_4_2 = uSystolicPE_300_io_randW_d;
  assign uSystolicPE_301_io_mac_done = mac_done_x_4[2];
  assign uSystolicPE_301_io_enable_i = enable_i_x_4[2];
  assign uSystolicPE_301_io_clear_i = clear_i_x_4[2];
  assign ifm_sign_x_4_3 = uSystolicPE_301_io_ifm_sign_d;
  assign ifm_dff_x_4_3 = uSystolicPE_301_io_ifm_dff_d;
  assign uSystolicPE_301_io_enable_w = enable_w_x_2[4];
  assign uSystolicPE_301_io_clear_w = clear_w_x_2[4];
  assign wght_sign_x_2_5 = uSystolicPE_301_io_wght_sign_d;
  assign wght_abs_x_2_5 = uSystolicPE_301_io_wght_abs_d;
  assign uSystolicPE_301_io_enable_o = enable_o_x_2[5];
  assign uSystolicPE_301_io_clear_o = clear_o_x_2[5];
  assign ofm_x_2_4 = uSystolicPE_301_io_ofm_d;
  assign randW_x_4_3 = uSystolicPE_301_io_randW_d;
  assign uSystolicPE_302_io_mac_done = mac_done_x_4[3];
  assign uSystolicPE_302_io_enable_i = enable_i_x_4[3];
  assign uSystolicPE_302_io_clear_i = clear_i_x_4[3];
  assign ifm_sign_x_4_4 = uSystolicPE_302_io_ifm_sign_d;
  assign ifm_dff_x_4_4 = uSystolicPE_302_io_ifm_dff_d;
  assign uSystolicPE_302_io_enable_w = enable_w_x_3[4];
  assign uSystolicPE_302_io_clear_w = clear_w_x_3[4];
  assign wght_sign_x_3_5 = uSystolicPE_302_io_wght_sign_d;
  assign wght_abs_x_3_5 = uSystolicPE_302_io_wght_abs_d;
  assign uSystolicPE_302_io_enable_o = enable_o_x_3[5];
  assign uSystolicPE_302_io_clear_o = clear_o_x_3[5];
  assign ofm_x_3_4 = uSystolicPE_302_io_ofm_d;
  assign randW_x_4_4 = uSystolicPE_302_io_randW_d;
  assign uSystolicPE_303_io_mac_done = mac_done_x_4[4];
  assign uSystolicPE_303_io_enable_i = enable_i_x_4[4];
  assign uSystolicPE_303_io_clear_i = clear_i_x_4[4];
  assign ifm_sign_x_4_5 = uSystolicPE_303_io_ifm_sign_d;
  assign ifm_dff_x_4_5 = uSystolicPE_303_io_ifm_dff_d;
  assign uSystolicPE_303_io_enable_w = enable_w_x_4[4];
  assign uSystolicPE_303_io_clear_w = clear_w_x_4[4];
  assign wght_sign_x_4_5 = uSystolicPE_303_io_wght_sign_d;
  assign wght_abs_x_4_5 = uSystolicPE_303_io_wght_abs_d;
  assign uSystolicPE_303_io_enable_o = enable_o_x_4[5];
  assign uSystolicPE_303_io_clear_o = clear_o_x_4[5];
  assign ofm_x_4_4 = uSystolicPE_303_io_ofm_d;
  assign randW_x_4_5 = uSystolicPE_303_io_randW_d;
  assign uSystolicPE_304_io_mac_done = mac_done_x_4[5];
  assign uSystolicPE_304_io_enable_i = enable_i_x_4[5];
  assign uSystolicPE_304_io_clear_i = clear_i_x_4[5];
  assign ifm_sign_x_4_6 = uSystolicPE_304_io_ifm_sign_d;
  assign ifm_dff_x_4_6 = uSystolicPE_304_io_ifm_dff_d;
  assign uSystolicPE_304_io_enable_w = enable_w_x_5[4];
  assign uSystolicPE_304_io_clear_w = clear_w_x_5[4];
  assign wght_sign_x_5_5 = uSystolicPE_304_io_wght_sign_d;
  assign wght_abs_x_5_5 = uSystolicPE_304_io_wght_abs_d;
  assign uSystolicPE_304_io_enable_o = enable_o_x_5[5];
  assign uSystolicPE_304_io_clear_o = clear_o_x_5[5];
  assign ofm_x_5_4 = uSystolicPE_304_io_ofm_d;
  assign randW_x_4_6 = uSystolicPE_304_io_randW_d;
  assign uSystolicPE_305_io_mac_done = mac_done_x_4[6];
  assign uSystolicPE_305_io_enable_i = enable_i_x_4[6];
  assign uSystolicPE_305_io_clear_i = clear_i_x_4[6];
  assign ifm_sign_x_4_7 = uSystolicPE_305_io_ifm_sign_d;
  assign ifm_dff_x_4_7 = uSystolicPE_305_io_ifm_dff_d;
  assign uSystolicPE_305_io_enable_w = enable_w_x_6[4];
  assign uSystolicPE_305_io_clear_w = clear_w_x_6[4];
  assign wght_sign_x_6_5 = uSystolicPE_305_io_wght_sign_d;
  assign wght_abs_x_6_5 = uSystolicPE_305_io_wght_abs_d;
  assign uSystolicPE_305_io_enable_o = enable_o_x_6[5];
  assign uSystolicPE_305_io_clear_o = clear_o_x_6[5];
  assign ofm_x_6_4 = uSystolicPE_305_io_ofm_d;
  assign randW_x_4_7 = uSystolicPE_305_io_randW_d;
  assign uSystolicPE_306_io_mac_done = mac_done_x_4[7];
  assign uSystolicPE_306_io_enable_i = enable_i_x_4[7];
  assign uSystolicPE_306_io_clear_i = clear_i_x_4[7];
  assign ifm_sign_x_4_8 = uSystolicPE_306_io_ifm_sign_d;
  assign ifm_dff_x_4_8 = uSystolicPE_306_io_ifm_dff_d;
  assign uSystolicPE_306_io_enable_w = enable_w_x_7[4];
  assign uSystolicPE_306_io_clear_w = clear_w_x_7[4];
  assign wght_sign_x_7_5 = uSystolicPE_306_io_wght_sign_d;
  assign wght_abs_x_7_5 = uSystolicPE_306_io_wght_abs_d;
  assign uSystolicPE_306_io_enable_o = enable_o_x_7[5];
  assign uSystolicPE_306_io_clear_o = clear_o_x_7[5];
  assign ofm_x_7_4 = uSystolicPE_306_io_ofm_d;
  assign randW_x_4_8 = uSystolicPE_306_io_randW_d;
  assign uSystolicPE_307_io_mac_done = mac_done_x_4[8];
  assign uSystolicPE_307_io_enable_i = enable_i_x_4[8];
  assign uSystolicPE_307_io_clear_i = clear_i_x_4[8];
  assign ifm_sign_x_4_9 = uSystolicPE_307_io_ifm_sign_d;
  assign ifm_dff_x_4_9 = uSystolicPE_307_io_ifm_dff_d;
  assign uSystolicPE_307_io_enable_w = enable_w_x_8[4];
  assign uSystolicPE_307_io_clear_w = clear_w_x_8[4];
  assign wght_sign_x_8_5 = uSystolicPE_307_io_wght_sign_d;
  assign wght_abs_x_8_5 = uSystolicPE_307_io_wght_abs_d;
  assign uSystolicPE_307_io_enable_o = enable_o_x_8[5];
  assign uSystolicPE_307_io_clear_o = clear_o_x_8[5];
  assign ofm_x_8_4 = uSystolicPE_307_io_ofm_d;
  assign randW_x_4_9 = uSystolicPE_307_io_randW_d;
  assign uSystolicPE_308_io_mac_done = mac_done_x_4[9];
  assign uSystolicPE_308_io_enable_i = enable_i_x_4[9];
  assign uSystolicPE_308_io_clear_i = clear_i_x_4[9];
  assign ifm_sign_x_4_10 = uSystolicPE_308_io_ifm_sign_d;
  assign ifm_dff_x_4_10 = uSystolicPE_308_io_ifm_dff_d;
  assign uSystolicPE_308_io_enable_w = enable_w_x_9[4];
  assign uSystolicPE_308_io_clear_w = clear_w_x_9[4];
  assign wght_sign_x_9_5 = uSystolicPE_308_io_wght_sign_d;
  assign wght_abs_x_9_5 = uSystolicPE_308_io_wght_abs_d;
  assign uSystolicPE_308_io_enable_o = enable_o_x_9[5];
  assign uSystolicPE_308_io_clear_o = clear_o_x_9[5];
  assign ofm_x_9_4 = uSystolicPE_308_io_ofm_d;
  assign randW_x_4_10 = uSystolicPE_308_io_randW_d;
  assign uSystolicPE_309_io_mac_done = mac_done_x_4[10];
  assign uSystolicPE_309_io_enable_i = enable_i_x_4[10];
  assign uSystolicPE_309_io_clear_i = clear_i_x_4[10];
  assign ifm_sign_x_4_11 = uSystolicPE_309_io_ifm_sign_d;
  assign ifm_dff_x_4_11 = uSystolicPE_309_io_ifm_dff_d;
  assign uSystolicPE_309_io_enable_w = enable_w_x_10[4];
  assign uSystolicPE_309_io_clear_w = clear_w_x_10[4];
  assign wght_sign_x_10_5 = uSystolicPE_309_io_wght_sign_d;
  assign wght_abs_x_10_5 = uSystolicPE_309_io_wght_abs_d;
  assign uSystolicPE_309_io_enable_o = enable_o_x_10[5];
  assign uSystolicPE_309_io_clear_o = clear_o_x_10[5];
  assign ofm_x_10_4 = uSystolicPE_309_io_ofm_d;
  assign randW_x_4_11 = uSystolicPE_309_io_randW_d;
  assign uSystolicPE_310_io_mac_done = mac_done_x_4[11];
  assign uSystolicPE_310_io_enable_i = enable_i_x_4[11];
  assign uSystolicPE_310_io_clear_i = clear_i_x_4[11];
  assign ifm_sign_x_4_12 = uSystolicPE_310_io_ifm_sign_d;
  assign ifm_dff_x_4_12 = uSystolicPE_310_io_ifm_dff_d;
  assign uSystolicPE_310_io_enable_w = enable_w_x_11[4];
  assign uSystolicPE_310_io_clear_w = clear_w_x_11[4];
  assign wght_sign_x_11_5 = uSystolicPE_310_io_wght_sign_d;
  assign wght_abs_x_11_5 = uSystolicPE_310_io_wght_abs_d;
  assign uSystolicPE_310_io_enable_o = enable_o_x_11[5];
  assign uSystolicPE_310_io_clear_o = clear_o_x_11[5];
  assign ofm_x_11_4 = uSystolicPE_310_io_ofm_d;
  assign randW_x_4_12 = uSystolicPE_310_io_randW_d;
  assign uSystolicPE_311_io_mac_done = mac_done_x_4[12];
  assign uSystolicPE_311_io_enable_i = enable_i_x_4[12];
  assign uSystolicPE_311_io_clear_i = clear_i_x_4[12];
  assign ifm_sign_x_4_13 = uSystolicPE_311_io_ifm_sign_d;
  assign ifm_dff_x_4_13 = uSystolicPE_311_io_ifm_dff_d;
  assign uSystolicPE_311_io_enable_w = enable_w_x_12[4];
  assign uSystolicPE_311_io_clear_w = clear_w_x_12[4];
  assign wght_sign_x_12_5 = uSystolicPE_311_io_wght_sign_d;
  assign wght_abs_x_12_5 = uSystolicPE_311_io_wght_abs_d;
  assign uSystolicPE_311_io_enable_o = enable_o_x_12[5];
  assign uSystolicPE_311_io_clear_o = clear_o_x_12[5];
  assign ofm_x_12_4 = uSystolicPE_311_io_ofm_d;
  assign randW_x_4_13 = uSystolicPE_311_io_randW_d;
  assign uSystolicPE_312_io_mac_done = mac_done_x_4[13];
  assign uSystolicPE_312_io_enable_i = enable_i_x_4[13];
  assign uSystolicPE_312_io_clear_i = clear_i_x_4[13];
  assign ifm_sign_x_4_14 = uSystolicPE_312_io_ifm_sign_d;
  assign ifm_dff_x_4_14 = uSystolicPE_312_io_ifm_dff_d;
  assign uSystolicPE_312_io_enable_w = enable_w_x_13[4];
  assign uSystolicPE_312_io_clear_w = clear_w_x_13[4];
  assign wght_sign_x_13_5 = uSystolicPE_312_io_wght_sign_d;
  assign wght_abs_x_13_5 = uSystolicPE_312_io_wght_abs_d;
  assign uSystolicPE_312_io_enable_o = enable_o_x_13[5];
  assign uSystolicPE_312_io_clear_o = clear_o_x_13[5];
  assign ofm_x_13_4 = uSystolicPE_312_io_ofm_d;
  assign randW_x_4_14 = uSystolicPE_312_io_randW_d;
  assign uSystolicPE_313_io_mac_done = mac_done_x_4[14];
  assign uSystolicPE_313_io_enable_i = enable_i_x_4[14];
  assign uSystolicPE_313_io_clear_i = clear_i_x_4[14];
  assign ifm_sign_x_4_15 = uSystolicPE_313_io_ifm_sign_d;
  assign ifm_dff_x_4_15 = uSystolicPE_313_io_ifm_dff_d;
  assign uSystolicPE_313_io_enable_w = enable_w_x_14[4];
  assign uSystolicPE_313_io_clear_w = clear_w_x_14[4];
  assign wght_sign_x_14_5 = uSystolicPE_313_io_wght_sign_d;
  assign wght_abs_x_14_5 = uSystolicPE_313_io_wght_abs_d;
  assign uSystolicPE_313_io_enable_o = enable_o_x_14[5];
  assign uSystolicPE_313_io_clear_o = clear_o_x_14[5];
  assign ofm_x_14_4 = uSystolicPE_313_io_ofm_d;
  assign randW_x_4_15 = uSystolicPE_313_io_randW_d;
  assign uSystolicPE_314_io_mac_done = mac_done_x_4[15];
  assign uSystolicPE_314_io_enable_i = enable_i_x_4[15];
  assign uSystolicPE_314_io_clear_i = clear_i_x_4[15];
  assign ifm_sign_x_4_16 = uSystolicPE_314_io_ifm_sign_d;
  assign ifm_dff_x_4_16 = uSystolicPE_314_io_ifm_dff_d;
  assign uSystolicPE_314_io_enable_w = enable_w_x_15[4];
  assign uSystolicPE_314_io_clear_w = clear_w_x_15[4];
  assign wght_sign_x_15_5 = uSystolicPE_314_io_wght_sign_d;
  assign wght_abs_x_15_5 = uSystolicPE_314_io_wght_abs_d;
  assign uSystolicPE_314_io_enable_o = enable_o_x_15[5];
  assign uSystolicPE_314_io_clear_o = clear_o_x_15[5];
  assign ofm_x_15_4 = uSystolicPE_314_io_ofm_d;
  assign randW_x_4_16 = uSystolicPE_314_io_randW_d;
  assign uSystolicPEBorder_21_io_mac_done = mac_done_x_5[0];
  assign uSystolicPEBorder_21_io_enable_i = enable_i_x_5[0];
  assign uSystolicPEBorder_21_io_clear_i = clear_i_x_5[0];
  assign ifm_sign_x_5_1 = uSystolicPEBorder_21_io_ifm_sign_d;
  assign ifm_dff_x_5_1 = uSystolicPEBorder_21_io_ifm_dff_d;
  assign uSystolicPEBorder_21_io_enable_w = enable_w_x_0[5];
  assign uSystolicPEBorder_21_io_clear_w = clear_w_x_0[5];
  assign wght_sign_x_0_6 = uSystolicPEBorder_21_io_wght_sign_d;
  assign wght_abs_x_0_6 = uSystolicPEBorder_21_io_wght_abs_d;
  assign uSystolicPEBorder_21_io_enable_o = enable_o_x_0[6];
  assign uSystolicPEBorder_21_io_clear_o = clear_o_x_0[6];
  assign ofm_x_0_5 = uSystolicPEBorder_21_io_ofm_d;
  assign randW_x_5_1 = uSystolicPEBorder_21_io_randW_d;
  assign uSystolicPE_315_io_mac_done = mac_done_x_5[1];
  assign uSystolicPE_315_io_enable_i = enable_i_x_5[1];
  assign uSystolicPE_315_io_clear_i = clear_i_x_5[1];
  assign ifm_sign_x_5_2 = uSystolicPE_315_io_ifm_sign_d;
  assign ifm_dff_x_5_2 = uSystolicPE_315_io_ifm_dff_d;
  assign uSystolicPE_315_io_enable_w = enable_w_x_1[5];
  assign uSystolicPE_315_io_clear_w = clear_w_x_1[5];
  assign wght_sign_x_1_6 = uSystolicPE_315_io_wght_sign_d;
  assign wght_abs_x_1_6 = uSystolicPE_315_io_wght_abs_d;
  assign uSystolicPE_315_io_enable_o = enable_o_x_1[6];
  assign uSystolicPE_315_io_clear_o = clear_o_x_1[6];
  assign ofm_x_1_5 = uSystolicPE_315_io_ofm_d;
  assign randW_x_5_2 = uSystolicPE_315_io_randW_d;
  assign uSystolicPE_316_io_mac_done = mac_done_x_5[2];
  assign uSystolicPE_316_io_enable_i = enable_i_x_5[2];
  assign uSystolicPE_316_io_clear_i = clear_i_x_5[2];
  assign ifm_sign_x_5_3 = uSystolicPE_316_io_ifm_sign_d;
  assign ifm_dff_x_5_3 = uSystolicPE_316_io_ifm_dff_d;
  assign uSystolicPE_316_io_enable_w = enable_w_x_2[5];
  assign uSystolicPE_316_io_clear_w = clear_w_x_2[5];
  assign wght_sign_x_2_6 = uSystolicPE_316_io_wght_sign_d;
  assign wght_abs_x_2_6 = uSystolicPE_316_io_wght_abs_d;
  assign uSystolicPE_316_io_enable_o = enable_o_x_2[6];
  assign uSystolicPE_316_io_clear_o = clear_o_x_2[6];
  assign ofm_x_2_5 = uSystolicPE_316_io_ofm_d;
  assign randW_x_5_3 = uSystolicPE_316_io_randW_d;
  assign uSystolicPE_317_io_mac_done = mac_done_x_5[3];
  assign uSystolicPE_317_io_enable_i = enable_i_x_5[3];
  assign uSystolicPE_317_io_clear_i = clear_i_x_5[3];
  assign ifm_sign_x_5_4 = uSystolicPE_317_io_ifm_sign_d;
  assign ifm_dff_x_5_4 = uSystolicPE_317_io_ifm_dff_d;
  assign uSystolicPE_317_io_enable_w = enable_w_x_3[5];
  assign uSystolicPE_317_io_clear_w = clear_w_x_3[5];
  assign wght_sign_x_3_6 = uSystolicPE_317_io_wght_sign_d;
  assign wght_abs_x_3_6 = uSystolicPE_317_io_wght_abs_d;
  assign uSystolicPE_317_io_enable_o = enable_o_x_3[6];
  assign uSystolicPE_317_io_clear_o = clear_o_x_3[6];
  assign ofm_x_3_5 = uSystolicPE_317_io_ofm_d;
  assign randW_x_5_4 = uSystolicPE_317_io_randW_d;
  assign uSystolicPE_318_io_mac_done = mac_done_x_5[4];
  assign uSystolicPE_318_io_enable_i = enable_i_x_5[4];
  assign uSystolicPE_318_io_clear_i = clear_i_x_5[4];
  assign ifm_sign_x_5_5 = uSystolicPE_318_io_ifm_sign_d;
  assign ifm_dff_x_5_5 = uSystolicPE_318_io_ifm_dff_d;
  assign uSystolicPE_318_io_enable_w = enable_w_x_4[5];
  assign uSystolicPE_318_io_clear_w = clear_w_x_4[5];
  assign wght_sign_x_4_6 = uSystolicPE_318_io_wght_sign_d;
  assign wght_abs_x_4_6 = uSystolicPE_318_io_wght_abs_d;
  assign uSystolicPE_318_io_enable_o = enable_o_x_4[6];
  assign uSystolicPE_318_io_clear_o = clear_o_x_4[6];
  assign ofm_x_4_5 = uSystolicPE_318_io_ofm_d;
  assign randW_x_5_5 = uSystolicPE_318_io_randW_d;
  assign uSystolicPE_319_io_mac_done = mac_done_x_5[5];
  assign uSystolicPE_319_io_enable_i = enable_i_x_5[5];
  assign uSystolicPE_319_io_clear_i = clear_i_x_5[5];
  assign ifm_sign_x_5_6 = uSystolicPE_319_io_ifm_sign_d;
  assign ifm_dff_x_5_6 = uSystolicPE_319_io_ifm_dff_d;
  assign uSystolicPE_319_io_enable_w = enable_w_x_5[5];
  assign uSystolicPE_319_io_clear_w = clear_w_x_5[5];
  assign wght_sign_x_5_6 = uSystolicPE_319_io_wght_sign_d;
  assign wght_abs_x_5_6 = uSystolicPE_319_io_wght_abs_d;
  assign uSystolicPE_319_io_enable_o = enable_o_x_5[6];
  assign uSystolicPE_319_io_clear_o = clear_o_x_5[6];
  assign ofm_x_5_5 = uSystolicPE_319_io_ofm_d;
  assign randW_x_5_6 = uSystolicPE_319_io_randW_d;
  assign uSystolicPE_320_io_mac_done = mac_done_x_5[6];
  assign uSystolicPE_320_io_enable_i = enable_i_x_5[6];
  assign uSystolicPE_320_io_clear_i = clear_i_x_5[6];
  assign ifm_sign_x_5_7 = uSystolicPE_320_io_ifm_sign_d;
  assign ifm_dff_x_5_7 = uSystolicPE_320_io_ifm_dff_d;
  assign uSystolicPE_320_io_enable_w = enable_w_x_6[5];
  assign uSystolicPE_320_io_clear_w = clear_w_x_6[5];
  assign wght_sign_x_6_6 = uSystolicPE_320_io_wght_sign_d;
  assign wght_abs_x_6_6 = uSystolicPE_320_io_wght_abs_d;
  assign uSystolicPE_320_io_enable_o = enable_o_x_6[6];
  assign uSystolicPE_320_io_clear_o = clear_o_x_6[6];
  assign ofm_x_6_5 = uSystolicPE_320_io_ofm_d;
  assign randW_x_5_7 = uSystolicPE_320_io_randW_d;
  assign uSystolicPE_321_io_mac_done = mac_done_x_5[7];
  assign uSystolicPE_321_io_enable_i = enable_i_x_5[7];
  assign uSystolicPE_321_io_clear_i = clear_i_x_5[7];
  assign ifm_sign_x_5_8 = uSystolicPE_321_io_ifm_sign_d;
  assign ifm_dff_x_5_8 = uSystolicPE_321_io_ifm_dff_d;
  assign uSystolicPE_321_io_enable_w = enable_w_x_7[5];
  assign uSystolicPE_321_io_clear_w = clear_w_x_7[5];
  assign wght_sign_x_7_6 = uSystolicPE_321_io_wght_sign_d;
  assign wght_abs_x_7_6 = uSystolicPE_321_io_wght_abs_d;
  assign uSystolicPE_321_io_enable_o = enable_o_x_7[6];
  assign uSystolicPE_321_io_clear_o = clear_o_x_7[6];
  assign ofm_x_7_5 = uSystolicPE_321_io_ofm_d;
  assign randW_x_5_8 = uSystolicPE_321_io_randW_d;
  assign uSystolicPE_322_io_mac_done = mac_done_x_5[8];
  assign uSystolicPE_322_io_enable_i = enable_i_x_5[8];
  assign uSystolicPE_322_io_clear_i = clear_i_x_5[8];
  assign ifm_sign_x_5_9 = uSystolicPE_322_io_ifm_sign_d;
  assign ifm_dff_x_5_9 = uSystolicPE_322_io_ifm_dff_d;
  assign uSystolicPE_322_io_enable_w = enable_w_x_8[5];
  assign uSystolicPE_322_io_clear_w = clear_w_x_8[5];
  assign wght_sign_x_8_6 = uSystolicPE_322_io_wght_sign_d;
  assign wght_abs_x_8_6 = uSystolicPE_322_io_wght_abs_d;
  assign uSystolicPE_322_io_enable_o = enable_o_x_8[6];
  assign uSystolicPE_322_io_clear_o = clear_o_x_8[6];
  assign ofm_x_8_5 = uSystolicPE_322_io_ofm_d;
  assign randW_x_5_9 = uSystolicPE_322_io_randW_d;
  assign uSystolicPE_323_io_mac_done = mac_done_x_5[9];
  assign uSystolicPE_323_io_enable_i = enable_i_x_5[9];
  assign uSystolicPE_323_io_clear_i = clear_i_x_5[9];
  assign ifm_sign_x_5_10 = uSystolicPE_323_io_ifm_sign_d;
  assign ifm_dff_x_5_10 = uSystolicPE_323_io_ifm_dff_d;
  assign uSystolicPE_323_io_enable_w = enable_w_x_9[5];
  assign uSystolicPE_323_io_clear_w = clear_w_x_9[5];
  assign wght_sign_x_9_6 = uSystolicPE_323_io_wght_sign_d;
  assign wght_abs_x_9_6 = uSystolicPE_323_io_wght_abs_d;
  assign uSystolicPE_323_io_enable_o = enable_o_x_9[6];
  assign uSystolicPE_323_io_clear_o = clear_o_x_9[6];
  assign ofm_x_9_5 = uSystolicPE_323_io_ofm_d;
  assign randW_x_5_10 = uSystolicPE_323_io_randW_d;
  assign uSystolicPE_324_io_mac_done = mac_done_x_5[10];
  assign uSystolicPE_324_io_enable_i = enable_i_x_5[10];
  assign uSystolicPE_324_io_clear_i = clear_i_x_5[10];
  assign ifm_sign_x_5_11 = uSystolicPE_324_io_ifm_sign_d;
  assign ifm_dff_x_5_11 = uSystolicPE_324_io_ifm_dff_d;
  assign uSystolicPE_324_io_enable_w = enable_w_x_10[5];
  assign uSystolicPE_324_io_clear_w = clear_w_x_10[5];
  assign wght_sign_x_10_6 = uSystolicPE_324_io_wght_sign_d;
  assign wght_abs_x_10_6 = uSystolicPE_324_io_wght_abs_d;
  assign uSystolicPE_324_io_enable_o = enable_o_x_10[6];
  assign uSystolicPE_324_io_clear_o = clear_o_x_10[6];
  assign ofm_x_10_5 = uSystolicPE_324_io_ofm_d;
  assign randW_x_5_11 = uSystolicPE_324_io_randW_d;
  assign uSystolicPE_325_io_mac_done = mac_done_x_5[11];
  assign uSystolicPE_325_io_enable_i = enable_i_x_5[11];
  assign uSystolicPE_325_io_clear_i = clear_i_x_5[11];
  assign ifm_sign_x_5_12 = uSystolicPE_325_io_ifm_sign_d;
  assign ifm_dff_x_5_12 = uSystolicPE_325_io_ifm_dff_d;
  assign uSystolicPE_325_io_enable_w = enable_w_x_11[5];
  assign uSystolicPE_325_io_clear_w = clear_w_x_11[5];
  assign wght_sign_x_11_6 = uSystolicPE_325_io_wght_sign_d;
  assign wght_abs_x_11_6 = uSystolicPE_325_io_wght_abs_d;
  assign uSystolicPE_325_io_enable_o = enable_o_x_11[6];
  assign uSystolicPE_325_io_clear_o = clear_o_x_11[6];
  assign ofm_x_11_5 = uSystolicPE_325_io_ofm_d;
  assign randW_x_5_12 = uSystolicPE_325_io_randW_d;
  assign uSystolicPE_326_io_mac_done = mac_done_x_5[12];
  assign uSystolicPE_326_io_enable_i = enable_i_x_5[12];
  assign uSystolicPE_326_io_clear_i = clear_i_x_5[12];
  assign ifm_sign_x_5_13 = uSystolicPE_326_io_ifm_sign_d;
  assign ifm_dff_x_5_13 = uSystolicPE_326_io_ifm_dff_d;
  assign uSystolicPE_326_io_enable_w = enable_w_x_12[5];
  assign uSystolicPE_326_io_clear_w = clear_w_x_12[5];
  assign wght_sign_x_12_6 = uSystolicPE_326_io_wght_sign_d;
  assign wght_abs_x_12_6 = uSystolicPE_326_io_wght_abs_d;
  assign uSystolicPE_326_io_enable_o = enable_o_x_12[6];
  assign uSystolicPE_326_io_clear_o = clear_o_x_12[6];
  assign ofm_x_12_5 = uSystolicPE_326_io_ofm_d;
  assign randW_x_5_13 = uSystolicPE_326_io_randW_d;
  assign uSystolicPE_327_io_mac_done = mac_done_x_5[13];
  assign uSystolicPE_327_io_enable_i = enable_i_x_5[13];
  assign uSystolicPE_327_io_clear_i = clear_i_x_5[13];
  assign ifm_sign_x_5_14 = uSystolicPE_327_io_ifm_sign_d;
  assign ifm_dff_x_5_14 = uSystolicPE_327_io_ifm_dff_d;
  assign uSystolicPE_327_io_enable_w = enable_w_x_13[5];
  assign uSystolicPE_327_io_clear_w = clear_w_x_13[5];
  assign wght_sign_x_13_6 = uSystolicPE_327_io_wght_sign_d;
  assign wght_abs_x_13_6 = uSystolicPE_327_io_wght_abs_d;
  assign uSystolicPE_327_io_enable_o = enable_o_x_13[6];
  assign uSystolicPE_327_io_clear_o = clear_o_x_13[6];
  assign ofm_x_13_5 = uSystolicPE_327_io_ofm_d;
  assign randW_x_5_14 = uSystolicPE_327_io_randW_d;
  assign uSystolicPE_328_io_mac_done = mac_done_x_5[14];
  assign uSystolicPE_328_io_enable_i = enable_i_x_5[14];
  assign uSystolicPE_328_io_clear_i = clear_i_x_5[14];
  assign ifm_sign_x_5_15 = uSystolicPE_328_io_ifm_sign_d;
  assign ifm_dff_x_5_15 = uSystolicPE_328_io_ifm_dff_d;
  assign uSystolicPE_328_io_enable_w = enable_w_x_14[5];
  assign uSystolicPE_328_io_clear_w = clear_w_x_14[5];
  assign wght_sign_x_14_6 = uSystolicPE_328_io_wght_sign_d;
  assign wght_abs_x_14_6 = uSystolicPE_328_io_wght_abs_d;
  assign uSystolicPE_328_io_enable_o = enable_o_x_14[6];
  assign uSystolicPE_328_io_clear_o = clear_o_x_14[6];
  assign ofm_x_14_5 = uSystolicPE_328_io_ofm_d;
  assign randW_x_5_15 = uSystolicPE_328_io_randW_d;
  assign uSystolicPE_329_io_mac_done = mac_done_x_5[15];
  assign uSystolicPE_329_io_enable_i = enable_i_x_5[15];
  assign uSystolicPE_329_io_clear_i = clear_i_x_5[15];
  assign ifm_sign_x_5_16 = uSystolicPE_329_io_ifm_sign_d;
  assign ifm_dff_x_5_16 = uSystolicPE_329_io_ifm_dff_d;
  assign uSystolicPE_329_io_enable_w = enable_w_x_15[5];
  assign uSystolicPE_329_io_clear_w = clear_w_x_15[5];
  assign wght_sign_x_15_6 = uSystolicPE_329_io_wght_sign_d;
  assign wght_abs_x_15_6 = uSystolicPE_329_io_wght_abs_d;
  assign uSystolicPE_329_io_enable_o = enable_o_x_15[6];
  assign uSystolicPE_329_io_clear_o = clear_o_x_15[6];
  assign ofm_x_15_5 = uSystolicPE_329_io_ofm_d;
  assign randW_x_5_16 = uSystolicPE_329_io_randW_d;
  assign uSystolicPEBorder_22_io_mac_done = mac_done_x_6[0];
  assign uSystolicPEBorder_22_io_enable_i = enable_i_x_6[0];
  assign uSystolicPEBorder_22_io_clear_i = clear_i_x_6[0];
  assign ifm_sign_x_6_1 = uSystolicPEBorder_22_io_ifm_sign_d;
  assign ifm_dff_x_6_1 = uSystolicPEBorder_22_io_ifm_dff_d;
  assign uSystolicPEBorder_22_io_enable_w = enable_w_x_0[6];
  assign uSystolicPEBorder_22_io_clear_w = clear_w_x_0[6];
  assign wght_sign_x_0_7 = uSystolicPEBorder_22_io_wght_sign_d;
  assign wght_abs_x_0_7 = uSystolicPEBorder_22_io_wght_abs_d;
  assign uSystolicPEBorder_22_io_enable_o = enable_o_x_0[7];
  assign uSystolicPEBorder_22_io_clear_o = clear_o_x_0[7];
  assign ofm_x_0_6 = uSystolicPEBorder_22_io_ofm_d;
  assign randW_x_6_1 = uSystolicPEBorder_22_io_randW_d;
  assign uSystolicPE_330_io_mac_done = mac_done_x_6[1];
  assign uSystolicPE_330_io_enable_i = enable_i_x_6[1];
  assign uSystolicPE_330_io_clear_i = clear_i_x_6[1];
  assign ifm_sign_x_6_2 = uSystolicPE_330_io_ifm_sign_d;
  assign ifm_dff_x_6_2 = uSystolicPE_330_io_ifm_dff_d;
  assign uSystolicPE_330_io_enable_w = enable_w_x_1[6];
  assign uSystolicPE_330_io_clear_w = clear_w_x_1[6];
  assign wght_sign_x_1_7 = uSystolicPE_330_io_wght_sign_d;
  assign wght_abs_x_1_7 = uSystolicPE_330_io_wght_abs_d;
  assign uSystolicPE_330_io_enable_o = enable_o_x_1[7];
  assign uSystolicPE_330_io_clear_o = clear_o_x_1[7];
  assign ofm_x_1_6 = uSystolicPE_330_io_ofm_d;
  assign randW_x_6_2 = uSystolicPE_330_io_randW_d;
  assign uSystolicPE_331_io_mac_done = mac_done_x_6[2];
  assign uSystolicPE_331_io_enable_i = enable_i_x_6[2];
  assign uSystolicPE_331_io_clear_i = clear_i_x_6[2];
  assign ifm_sign_x_6_3 = uSystolicPE_331_io_ifm_sign_d;
  assign ifm_dff_x_6_3 = uSystolicPE_331_io_ifm_dff_d;
  assign uSystolicPE_331_io_enable_w = enable_w_x_2[6];
  assign uSystolicPE_331_io_clear_w = clear_w_x_2[6];
  assign wght_sign_x_2_7 = uSystolicPE_331_io_wght_sign_d;
  assign wght_abs_x_2_7 = uSystolicPE_331_io_wght_abs_d;
  assign uSystolicPE_331_io_enable_o = enable_o_x_2[7];
  assign uSystolicPE_331_io_clear_o = clear_o_x_2[7];
  assign ofm_x_2_6 = uSystolicPE_331_io_ofm_d;
  assign randW_x_6_3 = uSystolicPE_331_io_randW_d;
  assign uSystolicPE_332_io_mac_done = mac_done_x_6[3];
  assign uSystolicPE_332_io_enable_i = enable_i_x_6[3];
  assign uSystolicPE_332_io_clear_i = clear_i_x_6[3];
  assign ifm_sign_x_6_4 = uSystolicPE_332_io_ifm_sign_d;
  assign ifm_dff_x_6_4 = uSystolicPE_332_io_ifm_dff_d;
  assign uSystolicPE_332_io_enable_w = enable_w_x_3[6];
  assign uSystolicPE_332_io_clear_w = clear_w_x_3[6];
  assign wght_sign_x_3_7 = uSystolicPE_332_io_wght_sign_d;
  assign wght_abs_x_3_7 = uSystolicPE_332_io_wght_abs_d;
  assign uSystolicPE_332_io_enable_o = enable_o_x_3[7];
  assign uSystolicPE_332_io_clear_o = clear_o_x_3[7];
  assign ofm_x_3_6 = uSystolicPE_332_io_ofm_d;
  assign randW_x_6_4 = uSystolicPE_332_io_randW_d;
  assign uSystolicPE_333_io_mac_done = mac_done_x_6[4];
  assign uSystolicPE_333_io_enable_i = enable_i_x_6[4];
  assign uSystolicPE_333_io_clear_i = clear_i_x_6[4];
  assign ifm_sign_x_6_5 = uSystolicPE_333_io_ifm_sign_d;
  assign ifm_dff_x_6_5 = uSystolicPE_333_io_ifm_dff_d;
  assign uSystolicPE_333_io_enable_w = enable_w_x_4[6];
  assign uSystolicPE_333_io_clear_w = clear_w_x_4[6];
  assign wght_sign_x_4_7 = uSystolicPE_333_io_wght_sign_d;
  assign wght_abs_x_4_7 = uSystolicPE_333_io_wght_abs_d;
  assign uSystolicPE_333_io_enable_o = enable_o_x_4[7];
  assign uSystolicPE_333_io_clear_o = clear_o_x_4[7];
  assign ofm_x_4_6 = uSystolicPE_333_io_ofm_d;
  assign randW_x_6_5 = uSystolicPE_333_io_randW_d;
  assign uSystolicPE_334_io_mac_done = mac_done_x_6[5];
  assign uSystolicPE_334_io_enable_i = enable_i_x_6[5];
  assign uSystolicPE_334_io_clear_i = clear_i_x_6[5];
  assign ifm_sign_x_6_6 = uSystolicPE_334_io_ifm_sign_d;
  assign ifm_dff_x_6_6 = uSystolicPE_334_io_ifm_dff_d;
  assign uSystolicPE_334_io_enable_w = enable_w_x_5[6];
  assign uSystolicPE_334_io_clear_w = clear_w_x_5[6];
  assign wght_sign_x_5_7 = uSystolicPE_334_io_wght_sign_d;
  assign wght_abs_x_5_7 = uSystolicPE_334_io_wght_abs_d;
  assign uSystolicPE_334_io_enable_o = enable_o_x_5[7];
  assign uSystolicPE_334_io_clear_o = clear_o_x_5[7];
  assign ofm_x_5_6 = uSystolicPE_334_io_ofm_d;
  assign randW_x_6_6 = uSystolicPE_334_io_randW_d;
  assign uSystolicPE_335_io_mac_done = mac_done_x_6[6];
  assign uSystolicPE_335_io_enable_i = enable_i_x_6[6];
  assign uSystolicPE_335_io_clear_i = clear_i_x_6[6];
  assign ifm_sign_x_6_7 = uSystolicPE_335_io_ifm_sign_d;
  assign ifm_dff_x_6_7 = uSystolicPE_335_io_ifm_dff_d;
  assign uSystolicPE_335_io_enable_w = enable_w_x_6[6];
  assign uSystolicPE_335_io_clear_w = clear_w_x_6[6];
  assign wght_sign_x_6_7 = uSystolicPE_335_io_wght_sign_d;
  assign wght_abs_x_6_7 = uSystolicPE_335_io_wght_abs_d;
  assign uSystolicPE_335_io_enable_o = enable_o_x_6[7];
  assign uSystolicPE_335_io_clear_o = clear_o_x_6[7];
  assign ofm_x_6_6 = uSystolicPE_335_io_ofm_d;
  assign randW_x_6_7 = uSystolicPE_335_io_randW_d;
  assign uSystolicPE_336_io_mac_done = mac_done_x_6[7];
  assign uSystolicPE_336_io_enable_i = enable_i_x_6[7];
  assign uSystolicPE_336_io_clear_i = clear_i_x_6[7];
  assign ifm_sign_x_6_8 = uSystolicPE_336_io_ifm_sign_d;
  assign ifm_dff_x_6_8 = uSystolicPE_336_io_ifm_dff_d;
  assign uSystolicPE_336_io_enable_w = enable_w_x_7[6];
  assign uSystolicPE_336_io_clear_w = clear_w_x_7[6];
  assign wght_sign_x_7_7 = uSystolicPE_336_io_wght_sign_d;
  assign wght_abs_x_7_7 = uSystolicPE_336_io_wght_abs_d;
  assign uSystolicPE_336_io_enable_o = enable_o_x_7[7];
  assign uSystolicPE_336_io_clear_o = clear_o_x_7[7];
  assign ofm_x_7_6 = uSystolicPE_336_io_ofm_d;
  assign randW_x_6_8 = uSystolicPE_336_io_randW_d;
  assign uSystolicPE_337_io_mac_done = mac_done_x_6[8];
  assign uSystolicPE_337_io_enable_i = enable_i_x_6[8];
  assign uSystolicPE_337_io_clear_i = clear_i_x_6[8];
  assign ifm_sign_x_6_9 = uSystolicPE_337_io_ifm_sign_d;
  assign ifm_dff_x_6_9 = uSystolicPE_337_io_ifm_dff_d;
  assign uSystolicPE_337_io_enable_w = enable_w_x_8[6];
  assign uSystolicPE_337_io_clear_w = clear_w_x_8[6];
  assign wght_sign_x_8_7 = uSystolicPE_337_io_wght_sign_d;
  assign wght_abs_x_8_7 = uSystolicPE_337_io_wght_abs_d;
  assign uSystolicPE_337_io_enable_o = enable_o_x_8[7];
  assign uSystolicPE_337_io_clear_o = clear_o_x_8[7];
  assign ofm_x_8_6 = uSystolicPE_337_io_ofm_d;
  assign randW_x_6_9 = uSystolicPE_337_io_randW_d;
  assign uSystolicPE_338_io_mac_done = mac_done_x_6[9];
  assign uSystolicPE_338_io_enable_i = enable_i_x_6[9];
  assign uSystolicPE_338_io_clear_i = clear_i_x_6[9];
  assign ifm_sign_x_6_10 = uSystolicPE_338_io_ifm_sign_d;
  assign ifm_dff_x_6_10 = uSystolicPE_338_io_ifm_dff_d;
  assign uSystolicPE_338_io_enable_w = enable_w_x_9[6];
  assign uSystolicPE_338_io_clear_w = clear_w_x_9[6];
  assign wght_sign_x_9_7 = uSystolicPE_338_io_wght_sign_d;
  assign wght_abs_x_9_7 = uSystolicPE_338_io_wght_abs_d;
  assign uSystolicPE_338_io_enable_o = enable_o_x_9[7];
  assign uSystolicPE_338_io_clear_o = clear_o_x_9[7];
  assign ofm_x_9_6 = uSystolicPE_338_io_ofm_d;
  assign randW_x_6_10 = uSystolicPE_338_io_randW_d;
  assign uSystolicPE_339_io_mac_done = mac_done_x_6[10];
  assign uSystolicPE_339_io_enable_i = enable_i_x_6[10];
  assign uSystolicPE_339_io_clear_i = clear_i_x_6[10];
  assign ifm_sign_x_6_11 = uSystolicPE_339_io_ifm_sign_d;
  assign ifm_dff_x_6_11 = uSystolicPE_339_io_ifm_dff_d;
  assign uSystolicPE_339_io_enable_w = enable_w_x_10[6];
  assign uSystolicPE_339_io_clear_w = clear_w_x_10[6];
  assign wght_sign_x_10_7 = uSystolicPE_339_io_wght_sign_d;
  assign wght_abs_x_10_7 = uSystolicPE_339_io_wght_abs_d;
  assign uSystolicPE_339_io_enable_o = enable_o_x_10[7];
  assign uSystolicPE_339_io_clear_o = clear_o_x_10[7];
  assign ofm_x_10_6 = uSystolicPE_339_io_ofm_d;
  assign randW_x_6_11 = uSystolicPE_339_io_randW_d;
  assign uSystolicPE_340_io_mac_done = mac_done_x_6[11];
  assign uSystolicPE_340_io_enable_i = enable_i_x_6[11];
  assign uSystolicPE_340_io_clear_i = clear_i_x_6[11];
  assign ifm_sign_x_6_12 = uSystolicPE_340_io_ifm_sign_d;
  assign ifm_dff_x_6_12 = uSystolicPE_340_io_ifm_dff_d;
  assign uSystolicPE_340_io_enable_w = enable_w_x_11[6];
  assign uSystolicPE_340_io_clear_w = clear_w_x_11[6];
  assign wght_sign_x_11_7 = uSystolicPE_340_io_wght_sign_d;
  assign wght_abs_x_11_7 = uSystolicPE_340_io_wght_abs_d;
  assign uSystolicPE_340_io_enable_o = enable_o_x_11[7];
  assign uSystolicPE_340_io_clear_o = clear_o_x_11[7];
  assign ofm_x_11_6 = uSystolicPE_340_io_ofm_d;
  assign randW_x_6_12 = uSystolicPE_340_io_randW_d;
  assign uSystolicPE_341_io_mac_done = mac_done_x_6[12];
  assign uSystolicPE_341_io_enable_i = enable_i_x_6[12];
  assign uSystolicPE_341_io_clear_i = clear_i_x_6[12];
  assign ifm_sign_x_6_13 = uSystolicPE_341_io_ifm_sign_d;
  assign ifm_dff_x_6_13 = uSystolicPE_341_io_ifm_dff_d;
  assign uSystolicPE_341_io_enable_w = enable_w_x_12[6];
  assign uSystolicPE_341_io_clear_w = clear_w_x_12[6];
  assign wght_sign_x_12_7 = uSystolicPE_341_io_wght_sign_d;
  assign wght_abs_x_12_7 = uSystolicPE_341_io_wght_abs_d;
  assign uSystolicPE_341_io_enable_o = enable_o_x_12[7];
  assign uSystolicPE_341_io_clear_o = clear_o_x_12[7];
  assign ofm_x_12_6 = uSystolicPE_341_io_ofm_d;
  assign randW_x_6_13 = uSystolicPE_341_io_randW_d;
  assign uSystolicPE_342_io_mac_done = mac_done_x_6[13];
  assign uSystolicPE_342_io_enable_i = enable_i_x_6[13];
  assign uSystolicPE_342_io_clear_i = clear_i_x_6[13];
  assign ifm_sign_x_6_14 = uSystolicPE_342_io_ifm_sign_d;
  assign ifm_dff_x_6_14 = uSystolicPE_342_io_ifm_dff_d;
  assign uSystolicPE_342_io_enable_w = enable_w_x_13[6];
  assign uSystolicPE_342_io_clear_w = clear_w_x_13[6];
  assign wght_sign_x_13_7 = uSystolicPE_342_io_wght_sign_d;
  assign wght_abs_x_13_7 = uSystolicPE_342_io_wght_abs_d;
  assign uSystolicPE_342_io_enable_o = enable_o_x_13[7];
  assign uSystolicPE_342_io_clear_o = clear_o_x_13[7];
  assign ofm_x_13_6 = uSystolicPE_342_io_ofm_d;
  assign randW_x_6_14 = uSystolicPE_342_io_randW_d;
  assign uSystolicPE_343_io_mac_done = mac_done_x_6[14];
  assign uSystolicPE_343_io_enable_i = enable_i_x_6[14];
  assign uSystolicPE_343_io_clear_i = clear_i_x_6[14];
  assign ifm_sign_x_6_15 = uSystolicPE_343_io_ifm_sign_d;
  assign ifm_dff_x_6_15 = uSystolicPE_343_io_ifm_dff_d;
  assign uSystolicPE_343_io_enable_w = enable_w_x_14[6];
  assign uSystolicPE_343_io_clear_w = clear_w_x_14[6];
  assign wght_sign_x_14_7 = uSystolicPE_343_io_wght_sign_d;
  assign wght_abs_x_14_7 = uSystolicPE_343_io_wght_abs_d;
  assign uSystolicPE_343_io_enable_o = enable_o_x_14[7];
  assign uSystolicPE_343_io_clear_o = clear_o_x_14[7];
  assign ofm_x_14_6 = uSystolicPE_343_io_ofm_d;
  assign randW_x_6_15 = uSystolicPE_343_io_randW_d;
  assign uSystolicPE_344_io_mac_done = mac_done_x_6[15];
  assign uSystolicPE_344_io_enable_i = enable_i_x_6[15];
  assign uSystolicPE_344_io_clear_i = clear_i_x_6[15];
  assign ifm_sign_x_6_16 = uSystolicPE_344_io_ifm_sign_d;
  assign ifm_dff_x_6_16 = uSystolicPE_344_io_ifm_dff_d;
  assign uSystolicPE_344_io_enable_w = enable_w_x_15[6];
  assign uSystolicPE_344_io_clear_w = clear_w_x_15[6];
  assign wght_sign_x_15_7 = uSystolicPE_344_io_wght_sign_d;
  assign wght_abs_x_15_7 = uSystolicPE_344_io_wght_abs_d;
  assign uSystolicPE_344_io_enable_o = enable_o_x_15[7];
  assign uSystolicPE_344_io_clear_o = clear_o_x_15[7];
  assign ofm_x_15_6 = uSystolicPE_344_io_ofm_d;
  assign randW_x_6_16 = uSystolicPE_344_io_randW_d;
  assign uSystolicPEBorder_23_io_mac_done = mac_done_x_7[0];
  assign uSystolicPEBorder_23_io_enable_i = enable_i_x_7[0];
  assign uSystolicPEBorder_23_io_clear_i = clear_i_x_7[0];
  assign ifm_sign_x_7_1 = uSystolicPEBorder_23_io_ifm_sign_d;
  assign ifm_dff_x_7_1 = uSystolicPEBorder_23_io_ifm_dff_d;
  assign uSystolicPEBorder_23_io_enable_w = enable_w_x_0[7];
  assign uSystolicPEBorder_23_io_clear_w = clear_w_x_0[7];
  assign wght_sign_x_0_8 = uSystolicPEBorder_23_io_wght_sign_d;
  assign wght_abs_x_0_8 = uSystolicPEBorder_23_io_wght_abs_d;
  assign uSystolicPEBorder_23_io_enable_o = enable_o_x_0[8];
  assign uSystolicPEBorder_23_io_clear_o = clear_o_x_0[8];
  assign ofm_x_0_7 = uSystolicPEBorder_23_io_ofm_d;
  assign randW_x_7_1 = uSystolicPEBorder_23_io_randW_d;
  assign uSystolicPE_345_io_mac_done = mac_done_x_7[1];
  assign uSystolicPE_345_io_enable_i = enable_i_x_7[1];
  assign uSystolicPE_345_io_clear_i = clear_i_x_7[1];
  assign ifm_sign_x_7_2 = uSystolicPE_345_io_ifm_sign_d;
  assign ifm_dff_x_7_2 = uSystolicPE_345_io_ifm_dff_d;
  assign uSystolicPE_345_io_enable_w = enable_w_x_1[7];
  assign uSystolicPE_345_io_clear_w = clear_w_x_1[7];
  assign wght_sign_x_1_8 = uSystolicPE_345_io_wght_sign_d;
  assign wght_abs_x_1_8 = uSystolicPE_345_io_wght_abs_d;
  assign uSystolicPE_345_io_enable_o = enable_o_x_1[8];
  assign uSystolicPE_345_io_clear_o = clear_o_x_1[8];
  assign ofm_x_1_7 = uSystolicPE_345_io_ofm_d;
  assign randW_x_7_2 = uSystolicPE_345_io_randW_d;
  assign uSystolicPE_346_io_mac_done = mac_done_x_7[2];
  assign uSystolicPE_346_io_enable_i = enable_i_x_7[2];
  assign uSystolicPE_346_io_clear_i = clear_i_x_7[2];
  assign ifm_sign_x_7_3 = uSystolicPE_346_io_ifm_sign_d;
  assign ifm_dff_x_7_3 = uSystolicPE_346_io_ifm_dff_d;
  assign uSystolicPE_346_io_enable_w = enable_w_x_2[7];
  assign uSystolicPE_346_io_clear_w = clear_w_x_2[7];
  assign wght_sign_x_2_8 = uSystolicPE_346_io_wght_sign_d;
  assign wght_abs_x_2_8 = uSystolicPE_346_io_wght_abs_d;
  assign uSystolicPE_346_io_enable_o = enable_o_x_2[8];
  assign uSystolicPE_346_io_clear_o = clear_o_x_2[8];
  assign ofm_x_2_7 = uSystolicPE_346_io_ofm_d;
  assign randW_x_7_3 = uSystolicPE_346_io_randW_d;
  assign uSystolicPE_347_io_mac_done = mac_done_x_7[3];
  assign uSystolicPE_347_io_enable_i = enable_i_x_7[3];
  assign uSystolicPE_347_io_clear_i = clear_i_x_7[3];
  assign ifm_sign_x_7_4 = uSystolicPE_347_io_ifm_sign_d;
  assign ifm_dff_x_7_4 = uSystolicPE_347_io_ifm_dff_d;
  assign uSystolicPE_347_io_enable_w = enable_w_x_3[7];
  assign uSystolicPE_347_io_clear_w = clear_w_x_3[7];
  assign wght_sign_x_3_8 = uSystolicPE_347_io_wght_sign_d;
  assign wght_abs_x_3_8 = uSystolicPE_347_io_wght_abs_d;
  assign uSystolicPE_347_io_enable_o = enable_o_x_3[8];
  assign uSystolicPE_347_io_clear_o = clear_o_x_3[8];
  assign ofm_x_3_7 = uSystolicPE_347_io_ofm_d;
  assign randW_x_7_4 = uSystolicPE_347_io_randW_d;
  assign uSystolicPE_348_io_mac_done = mac_done_x_7[4];
  assign uSystolicPE_348_io_enable_i = enable_i_x_7[4];
  assign uSystolicPE_348_io_clear_i = clear_i_x_7[4];
  assign ifm_sign_x_7_5 = uSystolicPE_348_io_ifm_sign_d;
  assign ifm_dff_x_7_5 = uSystolicPE_348_io_ifm_dff_d;
  assign uSystolicPE_348_io_enable_w = enable_w_x_4[7];
  assign uSystolicPE_348_io_clear_w = clear_w_x_4[7];
  assign wght_sign_x_4_8 = uSystolicPE_348_io_wght_sign_d;
  assign wght_abs_x_4_8 = uSystolicPE_348_io_wght_abs_d;
  assign uSystolicPE_348_io_enable_o = enable_o_x_4[8];
  assign uSystolicPE_348_io_clear_o = clear_o_x_4[8];
  assign ofm_x_4_7 = uSystolicPE_348_io_ofm_d;
  assign randW_x_7_5 = uSystolicPE_348_io_randW_d;
  assign uSystolicPE_349_io_mac_done = mac_done_x_7[5];
  assign uSystolicPE_349_io_enable_i = enable_i_x_7[5];
  assign uSystolicPE_349_io_clear_i = clear_i_x_7[5];
  assign ifm_sign_x_7_6 = uSystolicPE_349_io_ifm_sign_d;
  assign ifm_dff_x_7_6 = uSystolicPE_349_io_ifm_dff_d;
  assign uSystolicPE_349_io_enable_w = enable_w_x_5[7];
  assign uSystolicPE_349_io_clear_w = clear_w_x_5[7];
  assign wght_sign_x_5_8 = uSystolicPE_349_io_wght_sign_d;
  assign wght_abs_x_5_8 = uSystolicPE_349_io_wght_abs_d;
  assign uSystolicPE_349_io_enable_o = enable_o_x_5[8];
  assign uSystolicPE_349_io_clear_o = clear_o_x_5[8];
  assign ofm_x_5_7 = uSystolicPE_349_io_ofm_d;
  assign randW_x_7_6 = uSystolicPE_349_io_randW_d;
  assign uSystolicPE_350_io_mac_done = mac_done_x_7[6];
  assign uSystolicPE_350_io_enable_i = enable_i_x_7[6];
  assign uSystolicPE_350_io_clear_i = clear_i_x_7[6];
  assign ifm_sign_x_7_7 = uSystolicPE_350_io_ifm_sign_d;
  assign ifm_dff_x_7_7 = uSystolicPE_350_io_ifm_dff_d;
  assign uSystolicPE_350_io_enable_w = enable_w_x_6[7];
  assign uSystolicPE_350_io_clear_w = clear_w_x_6[7];
  assign wght_sign_x_6_8 = uSystolicPE_350_io_wght_sign_d;
  assign wght_abs_x_6_8 = uSystolicPE_350_io_wght_abs_d;
  assign uSystolicPE_350_io_enable_o = enable_o_x_6[8];
  assign uSystolicPE_350_io_clear_o = clear_o_x_6[8];
  assign ofm_x_6_7 = uSystolicPE_350_io_ofm_d;
  assign randW_x_7_7 = uSystolicPE_350_io_randW_d;
  assign uSystolicPE_351_io_mac_done = mac_done_x_7[7];
  assign uSystolicPE_351_io_enable_i = enable_i_x_7[7];
  assign uSystolicPE_351_io_clear_i = clear_i_x_7[7];
  assign ifm_sign_x_7_8 = uSystolicPE_351_io_ifm_sign_d;
  assign ifm_dff_x_7_8 = uSystolicPE_351_io_ifm_dff_d;
  assign uSystolicPE_351_io_enable_w = enable_w_x_7[7];
  assign uSystolicPE_351_io_clear_w = clear_w_x_7[7];
  assign wght_sign_x_7_8 = uSystolicPE_351_io_wght_sign_d;
  assign wght_abs_x_7_8 = uSystolicPE_351_io_wght_abs_d;
  assign uSystolicPE_351_io_enable_o = enable_o_x_7[8];
  assign uSystolicPE_351_io_clear_o = clear_o_x_7[8];
  assign ofm_x_7_7 = uSystolicPE_351_io_ofm_d;
  assign randW_x_7_8 = uSystolicPE_351_io_randW_d;
  assign uSystolicPE_352_io_mac_done = mac_done_x_7[8];
  assign uSystolicPE_352_io_enable_i = enable_i_x_7[8];
  assign uSystolicPE_352_io_clear_i = clear_i_x_7[8];
  assign ifm_sign_x_7_9 = uSystolicPE_352_io_ifm_sign_d;
  assign ifm_dff_x_7_9 = uSystolicPE_352_io_ifm_dff_d;
  assign uSystolicPE_352_io_enable_w = enable_w_x_8[7];
  assign uSystolicPE_352_io_clear_w = clear_w_x_8[7];
  assign wght_sign_x_8_8 = uSystolicPE_352_io_wght_sign_d;
  assign wght_abs_x_8_8 = uSystolicPE_352_io_wght_abs_d;
  assign uSystolicPE_352_io_enable_o = enable_o_x_8[8];
  assign uSystolicPE_352_io_clear_o = clear_o_x_8[8];
  assign ofm_x_8_7 = uSystolicPE_352_io_ofm_d;
  assign randW_x_7_9 = uSystolicPE_352_io_randW_d;
  assign uSystolicPE_353_io_mac_done = mac_done_x_7[9];
  assign uSystolicPE_353_io_enable_i = enable_i_x_7[9];
  assign uSystolicPE_353_io_clear_i = clear_i_x_7[9];
  assign ifm_sign_x_7_10 = uSystolicPE_353_io_ifm_sign_d;
  assign ifm_dff_x_7_10 = uSystolicPE_353_io_ifm_dff_d;
  assign uSystolicPE_353_io_enable_w = enable_w_x_9[7];
  assign uSystolicPE_353_io_clear_w = clear_w_x_9[7];
  assign wght_sign_x_9_8 = uSystolicPE_353_io_wght_sign_d;
  assign wght_abs_x_9_8 = uSystolicPE_353_io_wght_abs_d;
  assign uSystolicPE_353_io_enable_o = enable_o_x_9[8];
  assign uSystolicPE_353_io_clear_o = clear_o_x_9[8];
  assign ofm_x_9_7 = uSystolicPE_353_io_ofm_d;
  assign randW_x_7_10 = uSystolicPE_353_io_randW_d;
  assign uSystolicPE_354_io_mac_done = mac_done_x_7[10];
  assign uSystolicPE_354_io_enable_i = enable_i_x_7[10];
  assign uSystolicPE_354_io_clear_i = clear_i_x_7[10];
  assign ifm_sign_x_7_11 = uSystolicPE_354_io_ifm_sign_d;
  assign ifm_dff_x_7_11 = uSystolicPE_354_io_ifm_dff_d;
  assign uSystolicPE_354_io_enable_w = enable_w_x_10[7];
  assign uSystolicPE_354_io_clear_w = clear_w_x_10[7];
  assign wght_sign_x_10_8 = uSystolicPE_354_io_wght_sign_d;
  assign wght_abs_x_10_8 = uSystolicPE_354_io_wght_abs_d;
  assign uSystolicPE_354_io_enable_o = enable_o_x_10[8];
  assign uSystolicPE_354_io_clear_o = clear_o_x_10[8];
  assign ofm_x_10_7 = uSystolicPE_354_io_ofm_d;
  assign randW_x_7_11 = uSystolicPE_354_io_randW_d;
  assign uSystolicPE_355_io_mac_done = mac_done_x_7[11];
  assign uSystolicPE_355_io_enable_i = enable_i_x_7[11];
  assign uSystolicPE_355_io_clear_i = clear_i_x_7[11];
  assign ifm_sign_x_7_12 = uSystolicPE_355_io_ifm_sign_d;
  assign ifm_dff_x_7_12 = uSystolicPE_355_io_ifm_dff_d;
  assign uSystolicPE_355_io_enable_w = enable_w_x_11[7];
  assign uSystolicPE_355_io_clear_w = clear_w_x_11[7];
  assign wght_sign_x_11_8 = uSystolicPE_355_io_wght_sign_d;
  assign wght_abs_x_11_8 = uSystolicPE_355_io_wght_abs_d;
  assign uSystolicPE_355_io_enable_o = enable_o_x_11[8];
  assign uSystolicPE_355_io_clear_o = clear_o_x_11[8];
  assign ofm_x_11_7 = uSystolicPE_355_io_ofm_d;
  assign randW_x_7_12 = uSystolicPE_355_io_randW_d;
  assign uSystolicPE_356_io_mac_done = mac_done_x_7[12];
  assign uSystolicPE_356_io_enable_i = enable_i_x_7[12];
  assign uSystolicPE_356_io_clear_i = clear_i_x_7[12];
  assign ifm_sign_x_7_13 = uSystolicPE_356_io_ifm_sign_d;
  assign ifm_dff_x_7_13 = uSystolicPE_356_io_ifm_dff_d;
  assign uSystolicPE_356_io_enable_w = enable_w_x_12[7];
  assign uSystolicPE_356_io_clear_w = clear_w_x_12[7];
  assign wght_sign_x_12_8 = uSystolicPE_356_io_wght_sign_d;
  assign wght_abs_x_12_8 = uSystolicPE_356_io_wght_abs_d;
  assign uSystolicPE_356_io_enable_o = enable_o_x_12[8];
  assign uSystolicPE_356_io_clear_o = clear_o_x_12[8];
  assign ofm_x_12_7 = uSystolicPE_356_io_ofm_d;
  assign randW_x_7_13 = uSystolicPE_356_io_randW_d;
  assign uSystolicPE_357_io_mac_done = mac_done_x_7[13];
  assign uSystolicPE_357_io_enable_i = enable_i_x_7[13];
  assign uSystolicPE_357_io_clear_i = clear_i_x_7[13];
  assign ifm_sign_x_7_14 = uSystolicPE_357_io_ifm_sign_d;
  assign ifm_dff_x_7_14 = uSystolicPE_357_io_ifm_dff_d;
  assign uSystolicPE_357_io_enable_w = enable_w_x_13[7];
  assign uSystolicPE_357_io_clear_w = clear_w_x_13[7];
  assign wght_sign_x_13_8 = uSystolicPE_357_io_wght_sign_d;
  assign wght_abs_x_13_8 = uSystolicPE_357_io_wght_abs_d;
  assign uSystolicPE_357_io_enable_o = enable_o_x_13[8];
  assign uSystolicPE_357_io_clear_o = clear_o_x_13[8];
  assign ofm_x_13_7 = uSystolicPE_357_io_ofm_d;
  assign randW_x_7_14 = uSystolicPE_357_io_randW_d;
  assign uSystolicPE_358_io_mac_done = mac_done_x_7[14];
  assign uSystolicPE_358_io_enable_i = enable_i_x_7[14];
  assign uSystolicPE_358_io_clear_i = clear_i_x_7[14];
  assign ifm_sign_x_7_15 = uSystolicPE_358_io_ifm_sign_d;
  assign ifm_dff_x_7_15 = uSystolicPE_358_io_ifm_dff_d;
  assign uSystolicPE_358_io_enable_w = enable_w_x_14[7];
  assign uSystolicPE_358_io_clear_w = clear_w_x_14[7];
  assign wght_sign_x_14_8 = uSystolicPE_358_io_wght_sign_d;
  assign wght_abs_x_14_8 = uSystolicPE_358_io_wght_abs_d;
  assign uSystolicPE_358_io_enable_o = enable_o_x_14[8];
  assign uSystolicPE_358_io_clear_o = clear_o_x_14[8];
  assign ofm_x_14_7 = uSystolicPE_358_io_ofm_d;
  assign randW_x_7_15 = uSystolicPE_358_io_randW_d;
  assign uSystolicPE_359_io_mac_done = mac_done_x_7[15];
  assign uSystolicPE_359_io_enable_i = enable_i_x_7[15];
  assign uSystolicPE_359_io_clear_i = clear_i_x_7[15];
  assign ifm_sign_x_7_16 = uSystolicPE_359_io_ifm_sign_d;
  assign ifm_dff_x_7_16 = uSystolicPE_359_io_ifm_dff_d;
  assign uSystolicPE_359_io_enable_w = enable_w_x_15[7];
  assign uSystolicPE_359_io_clear_w = clear_w_x_15[7];
  assign wght_sign_x_15_8 = uSystolicPE_359_io_wght_sign_d;
  assign wght_abs_x_15_8 = uSystolicPE_359_io_wght_abs_d;
  assign uSystolicPE_359_io_enable_o = enable_o_x_15[8];
  assign uSystolicPE_359_io_clear_o = clear_o_x_15[8];
  assign ofm_x_15_7 = uSystolicPE_359_io_ofm_d;
  assign randW_x_7_16 = uSystolicPE_359_io_randW_d;
  assign uSystolicPEBorder_24_io_mac_done = mac_done_x_8[0];
  assign uSystolicPEBorder_24_io_enable_i = enable_i_x_8[0];
  assign uSystolicPEBorder_24_io_clear_i = clear_i_x_8[0];
  assign ifm_sign_x_8_1 = uSystolicPEBorder_24_io_ifm_sign_d;
  assign ifm_dff_x_8_1 = uSystolicPEBorder_24_io_ifm_dff_d;
  assign uSystolicPEBorder_24_io_enable_w = enable_w_x_0[8];
  assign uSystolicPEBorder_24_io_clear_w = clear_w_x_0[8];
  assign wght_sign_x_0_9 = uSystolicPEBorder_24_io_wght_sign_d;
  assign wght_abs_x_0_9 = uSystolicPEBorder_24_io_wght_abs_d;
  assign uSystolicPEBorder_24_io_enable_o = enable_o_x_0[9];
  assign uSystolicPEBorder_24_io_clear_o = clear_o_x_0[9];
  assign ofm_x_0_8 = uSystolicPEBorder_24_io_ofm_d;
  assign randW_x_8_1 = uSystolicPEBorder_24_io_randW_d;
  assign uSystolicPE_360_io_mac_done = mac_done_x_8[1];
  assign uSystolicPE_360_io_enable_i = enable_i_x_8[1];
  assign uSystolicPE_360_io_clear_i = clear_i_x_8[1];
  assign ifm_sign_x_8_2 = uSystolicPE_360_io_ifm_sign_d;
  assign ifm_dff_x_8_2 = uSystolicPE_360_io_ifm_dff_d;
  assign uSystolicPE_360_io_enable_w = enable_w_x_1[8];
  assign uSystolicPE_360_io_clear_w = clear_w_x_1[8];
  assign wght_sign_x_1_9 = uSystolicPE_360_io_wght_sign_d;
  assign wght_abs_x_1_9 = uSystolicPE_360_io_wght_abs_d;
  assign uSystolicPE_360_io_enable_o = enable_o_x_1[9];
  assign uSystolicPE_360_io_clear_o = clear_o_x_1[9];
  assign ofm_x_1_8 = uSystolicPE_360_io_ofm_d;
  assign randW_x_8_2 = uSystolicPE_360_io_randW_d;
  assign uSystolicPE_361_io_mac_done = mac_done_x_8[2];
  assign uSystolicPE_361_io_enable_i = enable_i_x_8[2];
  assign uSystolicPE_361_io_clear_i = clear_i_x_8[2];
  assign ifm_sign_x_8_3 = uSystolicPE_361_io_ifm_sign_d;
  assign ifm_dff_x_8_3 = uSystolicPE_361_io_ifm_dff_d;
  assign uSystolicPE_361_io_enable_w = enable_w_x_2[8];
  assign uSystolicPE_361_io_clear_w = clear_w_x_2[8];
  assign wght_sign_x_2_9 = uSystolicPE_361_io_wght_sign_d;
  assign wght_abs_x_2_9 = uSystolicPE_361_io_wght_abs_d;
  assign uSystolicPE_361_io_enable_o = enable_o_x_2[9];
  assign uSystolicPE_361_io_clear_o = clear_o_x_2[9];
  assign ofm_x_2_8 = uSystolicPE_361_io_ofm_d;
  assign randW_x_8_3 = uSystolicPE_361_io_randW_d;
  assign uSystolicPE_362_io_mac_done = mac_done_x_8[3];
  assign uSystolicPE_362_io_enable_i = enable_i_x_8[3];
  assign uSystolicPE_362_io_clear_i = clear_i_x_8[3];
  assign ifm_sign_x_8_4 = uSystolicPE_362_io_ifm_sign_d;
  assign ifm_dff_x_8_4 = uSystolicPE_362_io_ifm_dff_d;
  assign uSystolicPE_362_io_enable_w = enable_w_x_3[8];
  assign uSystolicPE_362_io_clear_w = clear_w_x_3[8];
  assign wght_sign_x_3_9 = uSystolicPE_362_io_wght_sign_d;
  assign wght_abs_x_3_9 = uSystolicPE_362_io_wght_abs_d;
  assign uSystolicPE_362_io_enable_o = enable_o_x_3[9];
  assign uSystolicPE_362_io_clear_o = clear_o_x_3[9];
  assign ofm_x_3_8 = uSystolicPE_362_io_ofm_d;
  assign randW_x_8_4 = uSystolicPE_362_io_randW_d;
  assign uSystolicPE_363_io_mac_done = mac_done_x_8[4];
  assign uSystolicPE_363_io_enable_i = enable_i_x_8[4];
  assign uSystolicPE_363_io_clear_i = clear_i_x_8[4];
  assign ifm_sign_x_8_5 = uSystolicPE_363_io_ifm_sign_d;
  assign ifm_dff_x_8_5 = uSystolicPE_363_io_ifm_dff_d;
  assign uSystolicPE_363_io_enable_w = enable_w_x_4[8];
  assign uSystolicPE_363_io_clear_w = clear_w_x_4[8];
  assign wght_sign_x_4_9 = uSystolicPE_363_io_wght_sign_d;
  assign wght_abs_x_4_9 = uSystolicPE_363_io_wght_abs_d;
  assign uSystolicPE_363_io_enable_o = enable_o_x_4[9];
  assign uSystolicPE_363_io_clear_o = clear_o_x_4[9];
  assign ofm_x_4_8 = uSystolicPE_363_io_ofm_d;
  assign randW_x_8_5 = uSystolicPE_363_io_randW_d;
  assign uSystolicPE_364_io_mac_done = mac_done_x_8[5];
  assign uSystolicPE_364_io_enable_i = enable_i_x_8[5];
  assign uSystolicPE_364_io_clear_i = clear_i_x_8[5];
  assign ifm_sign_x_8_6 = uSystolicPE_364_io_ifm_sign_d;
  assign ifm_dff_x_8_6 = uSystolicPE_364_io_ifm_dff_d;
  assign uSystolicPE_364_io_enable_w = enable_w_x_5[8];
  assign uSystolicPE_364_io_clear_w = clear_w_x_5[8];
  assign wght_sign_x_5_9 = uSystolicPE_364_io_wght_sign_d;
  assign wght_abs_x_5_9 = uSystolicPE_364_io_wght_abs_d;
  assign uSystolicPE_364_io_enable_o = enable_o_x_5[9];
  assign uSystolicPE_364_io_clear_o = clear_o_x_5[9];
  assign ofm_x_5_8 = uSystolicPE_364_io_ofm_d;
  assign randW_x_8_6 = uSystolicPE_364_io_randW_d;
  assign uSystolicPE_365_io_mac_done = mac_done_x_8[6];
  assign uSystolicPE_365_io_enable_i = enable_i_x_8[6];
  assign uSystolicPE_365_io_clear_i = clear_i_x_8[6];
  assign ifm_sign_x_8_7 = uSystolicPE_365_io_ifm_sign_d;
  assign ifm_dff_x_8_7 = uSystolicPE_365_io_ifm_dff_d;
  assign uSystolicPE_365_io_enable_w = enable_w_x_6[8];
  assign uSystolicPE_365_io_clear_w = clear_w_x_6[8];
  assign wght_sign_x_6_9 = uSystolicPE_365_io_wght_sign_d;
  assign wght_abs_x_6_9 = uSystolicPE_365_io_wght_abs_d;
  assign uSystolicPE_365_io_enable_o = enable_o_x_6[9];
  assign uSystolicPE_365_io_clear_o = clear_o_x_6[9];
  assign ofm_x_6_8 = uSystolicPE_365_io_ofm_d;
  assign randW_x_8_7 = uSystolicPE_365_io_randW_d;
  assign uSystolicPE_366_io_mac_done = mac_done_x_8[7];
  assign uSystolicPE_366_io_enable_i = enable_i_x_8[7];
  assign uSystolicPE_366_io_clear_i = clear_i_x_8[7];
  assign ifm_sign_x_8_8 = uSystolicPE_366_io_ifm_sign_d;
  assign ifm_dff_x_8_8 = uSystolicPE_366_io_ifm_dff_d;
  assign uSystolicPE_366_io_enable_w = enable_w_x_7[8];
  assign uSystolicPE_366_io_clear_w = clear_w_x_7[8];
  assign wght_sign_x_7_9 = uSystolicPE_366_io_wght_sign_d;
  assign wght_abs_x_7_9 = uSystolicPE_366_io_wght_abs_d;
  assign uSystolicPE_366_io_enable_o = enable_o_x_7[9];
  assign uSystolicPE_366_io_clear_o = clear_o_x_7[9];
  assign ofm_x_7_8 = uSystolicPE_366_io_ofm_d;
  assign randW_x_8_8 = uSystolicPE_366_io_randW_d;
  assign uSystolicPE_367_io_mac_done = mac_done_x_8[8];
  assign uSystolicPE_367_io_enable_i = enable_i_x_8[8];
  assign uSystolicPE_367_io_clear_i = clear_i_x_8[8];
  assign ifm_sign_x_8_9 = uSystolicPE_367_io_ifm_sign_d;
  assign ifm_dff_x_8_9 = uSystolicPE_367_io_ifm_dff_d;
  assign uSystolicPE_367_io_enable_w = enable_w_x_8[8];
  assign uSystolicPE_367_io_clear_w = clear_w_x_8[8];
  assign wght_sign_x_8_9 = uSystolicPE_367_io_wght_sign_d;
  assign wght_abs_x_8_9 = uSystolicPE_367_io_wght_abs_d;
  assign uSystolicPE_367_io_enable_o = enable_o_x_8[9];
  assign uSystolicPE_367_io_clear_o = clear_o_x_8[9];
  assign ofm_x_8_8 = uSystolicPE_367_io_ofm_d;
  assign randW_x_8_9 = uSystolicPE_367_io_randW_d;
  assign uSystolicPE_368_io_mac_done = mac_done_x_8[9];
  assign uSystolicPE_368_io_enable_i = enable_i_x_8[9];
  assign uSystolicPE_368_io_clear_i = clear_i_x_8[9];
  assign ifm_sign_x_8_10 = uSystolicPE_368_io_ifm_sign_d;
  assign ifm_dff_x_8_10 = uSystolicPE_368_io_ifm_dff_d;
  assign uSystolicPE_368_io_enable_w = enable_w_x_9[8];
  assign uSystolicPE_368_io_clear_w = clear_w_x_9[8];
  assign wght_sign_x_9_9 = uSystolicPE_368_io_wght_sign_d;
  assign wght_abs_x_9_9 = uSystolicPE_368_io_wght_abs_d;
  assign uSystolicPE_368_io_enable_o = enable_o_x_9[9];
  assign uSystolicPE_368_io_clear_o = clear_o_x_9[9];
  assign ofm_x_9_8 = uSystolicPE_368_io_ofm_d;
  assign randW_x_8_10 = uSystolicPE_368_io_randW_d;
  assign uSystolicPE_369_io_mac_done = mac_done_x_8[10];
  assign uSystolicPE_369_io_enable_i = enable_i_x_8[10];
  assign uSystolicPE_369_io_clear_i = clear_i_x_8[10];
  assign ifm_sign_x_8_11 = uSystolicPE_369_io_ifm_sign_d;
  assign ifm_dff_x_8_11 = uSystolicPE_369_io_ifm_dff_d;
  assign uSystolicPE_369_io_enable_w = enable_w_x_10[8];
  assign uSystolicPE_369_io_clear_w = clear_w_x_10[8];
  assign wght_sign_x_10_9 = uSystolicPE_369_io_wght_sign_d;
  assign wght_abs_x_10_9 = uSystolicPE_369_io_wght_abs_d;
  assign uSystolicPE_369_io_enable_o = enable_o_x_10[9];
  assign uSystolicPE_369_io_clear_o = clear_o_x_10[9];
  assign ofm_x_10_8 = uSystolicPE_369_io_ofm_d;
  assign randW_x_8_11 = uSystolicPE_369_io_randW_d;
  assign uSystolicPE_370_io_mac_done = mac_done_x_8[11];
  assign uSystolicPE_370_io_enable_i = enable_i_x_8[11];
  assign uSystolicPE_370_io_clear_i = clear_i_x_8[11];
  assign ifm_sign_x_8_12 = uSystolicPE_370_io_ifm_sign_d;
  assign ifm_dff_x_8_12 = uSystolicPE_370_io_ifm_dff_d;
  assign uSystolicPE_370_io_enable_w = enable_w_x_11[8];
  assign uSystolicPE_370_io_clear_w = clear_w_x_11[8];
  assign wght_sign_x_11_9 = uSystolicPE_370_io_wght_sign_d;
  assign wght_abs_x_11_9 = uSystolicPE_370_io_wght_abs_d;
  assign uSystolicPE_370_io_enable_o = enable_o_x_11[9];
  assign uSystolicPE_370_io_clear_o = clear_o_x_11[9];
  assign ofm_x_11_8 = uSystolicPE_370_io_ofm_d;
  assign randW_x_8_12 = uSystolicPE_370_io_randW_d;
  assign uSystolicPE_371_io_mac_done = mac_done_x_8[12];
  assign uSystolicPE_371_io_enable_i = enable_i_x_8[12];
  assign uSystolicPE_371_io_clear_i = clear_i_x_8[12];
  assign ifm_sign_x_8_13 = uSystolicPE_371_io_ifm_sign_d;
  assign ifm_dff_x_8_13 = uSystolicPE_371_io_ifm_dff_d;
  assign uSystolicPE_371_io_enable_w = enable_w_x_12[8];
  assign uSystolicPE_371_io_clear_w = clear_w_x_12[8];
  assign wght_sign_x_12_9 = uSystolicPE_371_io_wght_sign_d;
  assign wght_abs_x_12_9 = uSystolicPE_371_io_wght_abs_d;
  assign uSystolicPE_371_io_enable_o = enable_o_x_12[9];
  assign uSystolicPE_371_io_clear_o = clear_o_x_12[9];
  assign ofm_x_12_8 = uSystolicPE_371_io_ofm_d;
  assign randW_x_8_13 = uSystolicPE_371_io_randW_d;
  assign uSystolicPE_372_io_mac_done = mac_done_x_8[13];
  assign uSystolicPE_372_io_enable_i = enable_i_x_8[13];
  assign uSystolicPE_372_io_clear_i = clear_i_x_8[13];
  assign ifm_sign_x_8_14 = uSystolicPE_372_io_ifm_sign_d;
  assign ifm_dff_x_8_14 = uSystolicPE_372_io_ifm_dff_d;
  assign uSystolicPE_372_io_enable_w = enable_w_x_13[8];
  assign uSystolicPE_372_io_clear_w = clear_w_x_13[8];
  assign wght_sign_x_13_9 = uSystolicPE_372_io_wght_sign_d;
  assign wght_abs_x_13_9 = uSystolicPE_372_io_wght_abs_d;
  assign uSystolicPE_372_io_enable_o = enable_o_x_13[9];
  assign uSystolicPE_372_io_clear_o = clear_o_x_13[9];
  assign ofm_x_13_8 = uSystolicPE_372_io_ofm_d;
  assign randW_x_8_14 = uSystolicPE_372_io_randW_d;
  assign uSystolicPE_373_io_mac_done = mac_done_x_8[14];
  assign uSystolicPE_373_io_enable_i = enable_i_x_8[14];
  assign uSystolicPE_373_io_clear_i = clear_i_x_8[14];
  assign ifm_sign_x_8_15 = uSystolicPE_373_io_ifm_sign_d;
  assign ifm_dff_x_8_15 = uSystolicPE_373_io_ifm_dff_d;
  assign uSystolicPE_373_io_enable_w = enable_w_x_14[8];
  assign uSystolicPE_373_io_clear_w = clear_w_x_14[8];
  assign wght_sign_x_14_9 = uSystolicPE_373_io_wght_sign_d;
  assign wght_abs_x_14_9 = uSystolicPE_373_io_wght_abs_d;
  assign uSystolicPE_373_io_enable_o = enable_o_x_14[9];
  assign uSystolicPE_373_io_clear_o = clear_o_x_14[9];
  assign ofm_x_14_8 = uSystolicPE_373_io_ofm_d;
  assign randW_x_8_15 = uSystolicPE_373_io_randW_d;
  assign uSystolicPE_374_io_mac_done = mac_done_x_8[15];
  assign uSystolicPE_374_io_enable_i = enable_i_x_8[15];
  assign uSystolicPE_374_io_clear_i = clear_i_x_8[15];
  assign ifm_sign_x_8_16 = uSystolicPE_374_io_ifm_sign_d;
  assign ifm_dff_x_8_16 = uSystolicPE_374_io_ifm_dff_d;
  assign uSystolicPE_374_io_enable_w = enable_w_x_15[8];
  assign uSystolicPE_374_io_clear_w = clear_w_x_15[8];
  assign wght_sign_x_15_9 = uSystolicPE_374_io_wght_sign_d;
  assign wght_abs_x_15_9 = uSystolicPE_374_io_wght_abs_d;
  assign uSystolicPE_374_io_enable_o = enable_o_x_15[9];
  assign uSystolicPE_374_io_clear_o = clear_o_x_15[9];
  assign ofm_x_15_8 = uSystolicPE_374_io_ofm_d;
  assign randW_x_8_16 = uSystolicPE_374_io_randW_d;
  assign uSystolicPEBorder_25_io_mac_done = mac_done_x_9[0];
  assign uSystolicPEBorder_25_io_enable_i = enable_i_x_9[0];
  assign uSystolicPEBorder_25_io_clear_i = clear_i_x_9[0];
  assign ifm_sign_x_9_1 = uSystolicPEBorder_25_io_ifm_sign_d;
  assign ifm_dff_x_9_1 = uSystolicPEBorder_25_io_ifm_dff_d;
  assign uSystolicPEBorder_25_io_enable_w = enable_w_x_0[9];
  assign uSystolicPEBorder_25_io_clear_w = clear_w_x_0[9];
  assign wght_sign_x_0_10 = uSystolicPEBorder_25_io_wght_sign_d;
  assign wght_abs_x_0_10 = uSystolicPEBorder_25_io_wght_abs_d;
  assign uSystolicPEBorder_25_io_enable_o = enable_o_x_0[10];
  assign uSystolicPEBorder_25_io_clear_o = clear_o_x_0[10];
  assign ofm_x_0_9 = uSystolicPEBorder_25_io_ofm_d;
  assign randW_x_9_1 = uSystolicPEBorder_25_io_randW_d;
  assign uSystolicPE_375_io_mac_done = mac_done_x_9[1];
  assign uSystolicPE_375_io_enable_i = enable_i_x_9[1];
  assign uSystolicPE_375_io_clear_i = clear_i_x_9[1];
  assign ifm_sign_x_9_2 = uSystolicPE_375_io_ifm_sign_d;
  assign ifm_dff_x_9_2 = uSystolicPE_375_io_ifm_dff_d;
  assign uSystolicPE_375_io_enable_w = enable_w_x_1[9];
  assign uSystolicPE_375_io_clear_w = clear_w_x_1[9];
  assign wght_sign_x_1_10 = uSystolicPE_375_io_wght_sign_d;
  assign wght_abs_x_1_10 = uSystolicPE_375_io_wght_abs_d;
  assign uSystolicPE_375_io_enable_o = enable_o_x_1[10];
  assign uSystolicPE_375_io_clear_o = clear_o_x_1[10];
  assign ofm_x_1_9 = uSystolicPE_375_io_ofm_d;
  assign randW_x_9_2 = uSystolicPE_375_io_randW_d;
  assign uSystolicPE_376_io_mac_done = mac_done_x_9[2];
  assign uSystolicPE_376_io_enable_i = enable_i_x_9[2];
  assign uSystolicPE_376_io_clear_i = clear_i_x_9[2];
  assign ifm_sign_x_9_3 = uSystolicPE_376_io_ifm_sign_d;
  assign ifm_dff_x_9_3 = uSystolicPE_376_io_ifm_dff_d;
  assign uSystolicPE_376_io_enable_w = enable_w_x_2[9];
  assign uSystolicPE_376_io_clear_w = clear_w_x_2[9];
  assign wght_sign_x_2_10 = uSystolicPE_376_io_wght_sign_d;
  assign wght_abs_x_2_10 = uSystolicPE_376_io_wght_abs_d;
  assign uSystolicPE_376_io_enable_o = enable_o_x_2[10];
  assign uSystolicPE_376_io_clear_o = clear_o_x_2[10];
  assign ofm_x_2_9 = uSystolicPE_376_io_ofm_d;
  assign randW_x_9_3 = uSystolicPE_376_io_randW_d;
  assign uSystolicPE_377_io_mac_done = mac_done_x_9[3];
  assign uSystolicPE_377_io_enable_i = enable_i_x_9[3];
  assign uSystolicPE_377_io_clear_i = clear_i_x_9[3];
  assign ifm_sign_x_9_4 = uSystolicPE_377_io_ifm_sign_d;
  assign ifm_dff_x_9_4 = uSystolicPE_377_io_ifm_dff_d;
  assign uSystolicPE_377_io_enable_w = enable_w_x_3[9];
  assign uSystolicPE_377_io_clear_w = clear_w_x_3[9];
  assign wght_sign_x_3_10 = uSystolicPE_377_io_wght_sign_d;
  assign wght_abs_x_3_10 = uSystolicPE_377_io_wght_abs_d;
  assign uSystolicPE_377_io_enable_o = enable_o_x_3[10];
  assign uSystolicPE_377_io_clear_o = clear_o_x_3[10];
  assign ofm_x_3_9 = uSystolicPE_377_io_ofm_d;
  assign randW_x_9_4 = uSystolicPE_377_io_randW_d;
  assign uSystolicPE_378_io_mac_done = mac_done_x_9[4];
  assign uSystolicPE_378_io_enable_i = enable_i_x_9[4];
  assign uSystolicPE_378_io_clear_i = clear_i_x_9[4];
  assign ifm_sign_x_9_5 = uSystolicPE_378_io_ifm_sign_d;
  assign ifm_dff_x_9_5 = uSystolicPE_378_io_ifm_dff_d;
  assign uSystolicPE_378_io_enable_w = enable_w_x_4[9];
  assign uSystolicPE_378_io_clear_w = clear_w_x_4[9];
  assign wght_sign_x_4_10 = uSystolicPE_378_io_wght_sign_d;
  assign wght_abs_x_4_10 = uSystolicPE_378_io_wght_abs_d;
  assign uSystolicPE_378_io_enable_o = enable_o_x_4[10];
  assign uSystolicPE_378_io_clear_o = clear_o_x_4[10];
  assign ofm_x_4_9 = uSystolicPE_378_io_ofm_d;
  assign randW_x_9_5 = uSystolicPE_378_io_randW_d;
  assign uSystolicPE_379_io_mac_done = mac_done_x_9[5];
  assign uSystolicPE_379_io_enable_i = enable_i_x_9[5];
  assign uSystolicPE_379_io_clear_i = clear_i_x_9[5];
  assign ifm_sign_x_9_6 = uSystolicPE_379_io_ifm_sign_d;
  assign ifm_dff_x_9_6 = uSystolicPE_379_io_ifm_dff_d;
  assign uSystolicPE_379_io_enable_w = enable_w_x_5[9];
  assign uSystolicPE_379_io_clear_w = clear_w_x_5[9];
  assign wght_sign_x_5_10 = uSystolicPE_379_io_wght_sign_d;
  assign wght_abs_x_5_10 = uSystolicPE_379_io_wght_abs_d;
  assign uSystolicPE_379_io_enable_o = enable_o_x_5[10];
  assign uSystolicPE_379_io_clear_o = clear_o_x_5[10];
  assign ofm_x_5_9 = uSystolicPE_379_io_ofm_d;
  assign randW_x_9_6 = uSystolicPE_379_io_randW_d;
  assign uSystolicPE_380_io_mac_done = mac_done_x_9[6];
  assign uSystolicPE_380_io_enable_i = enable_i_x_9[6];
  assign uSystolicPE_380_io_clear_i = clear_i_x_9[6];
  assign ifm_sign_x_9_7 = uSystolicPE_380_io_ifm_sign_d;
  assign ifm_dff_x_9_7 = uSystolicPE_380_io_ifm_dff_d;
  assign uSystolicPE_380_io_enable_w = enable_w_x_6[9];
  assign uSystolicPE_380_io_clear_w = clear_w_x_6[9];
  assign wght_sign_x_6_10 = uSystolicPE_380_io_wght_sign_d;
  assign wght_abs_x_6_10 = uSystolicPE_380_io_wght_abs_d;
  assign uSystolicPE_380_io_enable_o = enable_o_x_6[10];
  assign uSystolicPE_380_io_clear_o = clear_o_x_6[10];
  assign ofm_x_6_9 = uSystolicPE_380_io_ofm_d;
  assign randW_x_9_7 = uSystolicPE_380_io_randW_d;
  assign uSystolicPE_381_io_mac_done = mac_done_x_9[7];
  assign uSystolicPE_381_io_enable_i = enable_i_x_9[7];
  assign uSystolicPE_381_io_clear_i = clear_i_x_9[7];
  assign ifm_sign_x_9_8 = uSystolicPE_381_io_ifm_sign_d;
  assign ifm_dff_x_9_8 = uSystolicPE_381_io_ifm_dff_d;
  assign uSystolicPE_381_io_enable_w = enable_w_x_7[9];
  assign uSystolicPE_381_io_clear_w = clear_w_x_7[9];
  assign wght_sign_x_7_10 = uSystolicPE_381_io_wght_sign_d;
  assign wght_abs_x_7_10 = uSystolicPE_381_io_wght_abs_d;
  assign uSystolicPE_381_io_enable_o = enable_o_x_7[10];
  assign uSystolicPE_381_io_clear_o = clear_o_x_7[10];
  assign ofm_x_7_9 = uSystolicPE_381_io_ofm_d;
  assign randW_x_9_8 = uSystolicPE_381_io_randW_d;
  assign uSystolicPE_382_io_mac_done = mac_done_x_9[8];
  assign uSystolicPE_382_io_enable_i = enable_i_x_9[8];
  assign uSystolicPE_382_io_clear_i = clear_i_x_9[8];
  assign ifm_sign_x_9_9 = uSystolicPE_382_io_ifm_sign_d;
  assign ifm_dff_x_9_9 = uSystolicPE_382_io_ifm_dff_d;
  assign uSystolicPE_382_io_enable_w = enable_w_x_8[9];
  assign uSystolicPE_382_io_clear_w = clear_w_x_8[9];
  assign wght_sign_x_8_10 = uSystolicPE_382_io_wght_sign_d;
  assign wght_abs_x_8_10 = uSystolicPE_382_io_wght_abs_d;
  assign uSystolicPE_382_io_enable_o = enable_o_x_8[10];
  assign uSystolicPE_382_io_clear_o = clear_o_x_8[10];
  assign ofm_x_8_9 = uSystolicPE_382_io_ofm_d;
  assign randW_x_9_9 = uSystolicPE_382_io_randW_d;
  assign uSystolicPE_383_io_mac_done = mac_done_x_9[9];
  assign uSystolicPE_383_io_enable_i = enable_i_x_9[9];
  assign uSystolicPE_383_io_clear_i = clear_i_x_9[9];
  assign ifm_sign_x_9_10 = uSystolicPE_383_io_ifm_sign_d;
  assign ifm_dff_x_9_10 = uSystolicPE_383_io_ifm_dff_d;
  assign uSystolicPE_383_io_enable_w = enable_w_x_9[9];
  assign uSystolicPE_383_io_clear_w = clear_w_x_9[9];
  assign wght_sign_x_9_10 = uSystolicPE_383_io_wght_sign_d;
  assign wght_abs_x_9_10 = uSystolicPE_383_io_wght_abs_d;
  assign uSystolicPE_383_io_enable_o = enable_o_x_9[10];
  assign uSystolicPE_383_io_clear_o = clear_o_x_9[10];
  assign ofm_x_9_9 = uSystolicPE_383_io_ofm_d;
  assign randW_x_9_10 = uSystolicPE_383_io_randW_d;
  assign uSystolicPE_384_io_mac_done = mac_done_x_9[10];
  assign uSystolicPE_384_io_enable_i = enable_i_x_9[10];
  assign uSystolicPE_384_io_clear_i = clear_i_x_9[10];
  assign ifm_sign_x_9_11 = uSystolicPE_384_io_ifm_sign_d;
  assign ifm_dff_x_9_11 = uSystolicPE_384_io_ifm_dff_d;
  assign uSystolicPE_384_io_enable_w = enable_w_x_10[9];
  assign uSystolicPE_384_io_clear_w = clear_w_x_10[9];
  assign wght_sign_x_10_10 = uSystolicPE_384_io_wght_sign_d;
  assign wght_abs_x_10_10 = uSystolicPE_384_io_wght_abs_d;
  assign uSystolicPE_384_io_enable_o = enable_o_x_10[10];
  assign uSystolicPE_384_io_clear_o = clear_o_x_10[10];
  assign ofm_x_10_9 = uSystolicPE_384_io_ofm_d;
  assign randW_x_9_11 = uSystolicPE_384_io_randW_d;
  assign uSystolicPE_385_io_mac_done = mac_done_x_9[11];
  assign uSystolicPE_385_io_enable_i = enable_i_x_9[11];
  assign uSystolicPE_385_io_clear_i = clear_i_x_9[11];
  assign ifm_sign_x_9_12 = uSystolicPE_385_io_ifm_sign_d;
  assign ifm_dff_x_9_12 = uSystolicPE_385_io_ifm_dff_d;
  assign uSystolicPE_385_io_enable_w = enable_w_x_11[9];
  assign uSystolicPE_385_io_clear_w = clear_w_x_11[9];
  assign wght_sign_x_11_10 = uSystolicPE_385_io_wght_sign_d;
  assign wght_abs_x_11_10 = uSystolicPE_385_io_wght_abs_d;
  assign uSystolicPE_385_io_enable_o = enable_o_x_11[10];
  assign uSystolicPE_385_io_clear_o = clear_o_x_11[10];
  assign ofm_x_11_9 = uSystolicPE_385_io_ofm_d;
  assign randW_x_9_12 = uSystolicPE_385_io_randW_d;
  assign uSystolicPE_386_io_mac_done = mac_done_x_9[12];
  assign uSystolicPE_386_io_enable_i = enable_i_x_9[12];
  assign uSystolicPE_386_io_clear_i = clear_i_x_9[12];
  assign ifm_sign_x_9_13 = uSystolicPE_386_io_ifm_sign_d;
  assign ifm_dff_x_9_13 = uSystolicPE_386_io_ifm_dff_d;
  assign uSystolicPE_386_io_enable_w = enable_w_x_12[9];
  assign uSystolicPE_386_io_clear_w = clear_w_x_12[9];
  assign wght_sign_x_12_10 = uSystolicPE_386_io_wght_sign_d;
  assign wght_abs_x_12_10 = uSystolicPE_386_io_wght_abs_d;
  assign uSystolicPE_386_io_enable_o = enable_o_x_12[10];
  assign uSystolicPE_386_io_clear_o = clear_o_x_12[10];
  assign ofm_x_12_9 = uSystolicPE_386_io_ofm_d;
  assign randW_x_9_13 = uSystolicPE_386_io_randW_d;
  assign uSystolicPE_387_io_mac_done = mac_done_x_9[13];
  assign uSystolicPE_387_io_enable_i = enable_i_x_9[13];
  assign uSystolicPE_387_io_clear_i = clear_i_x_9[13];
  assign ifm_sign_x_9_14 = uSystolicPE_387_io_ifm_sign_d;
  assign ifm_dff_x_9_14 = uSystolicPE_387_io_ifm_dff_d;
  assign uSystolicPE_387_io_enable_w = enable_w_x_13[9];
  assign uSystolicPE_387_io_clear_w = clear_w_x_13[9];
  assign wght_sign_x_13_10 = uSystolicPE_387_io_wght_sign_d;
  assign wght_abs_x_13_10 = uSystolicPE_387_io_wght_abs_d;
  assign uSystolicPE_387_io_enable_o = enable_o_x_13[10];
  assign uSystolicPE_387_io_clear_o = clear_o_x_13[10];
  assign ofm_x_13_9 = uSystolicPE_387_io_ofm_d;
  assign randW_x_9_14 = uSystolicPE_387_io_randW_d;
  assign uSystolicPE_388_io_mac_done = mac_done_x_9[14];
  assign uSystolicPE_388_io_enable_i = enable_i_x_9[14];
  assign uSystolicPE_388_io_clear_i = clear_i_x_9[14];
  assign ifm_sign_x_9_15 = uSystolicPE_388_io_ifm_sign_d;
  assign ifm_dff_x_9_15 = uSystolicPE_388_io_ifm_dff_d;
  assign uSystolicPE_388_io_enable_w = enable_w_x_14[9];
  assign uSystolicPE_388_io_clear_w = clear_w_x_14[9];
  assign wght_sign_x_14_10 = uSystolicPE_388_io_wght_sign_d;
  assign wght_abs_x_14_10 = uSystolicPE_388_io_wght_abs_d;
  assign uSystolicPE_388_io_enable_o = enable_o_x_14[10];
  assign uSystolicPE_388_io_clear_o = clear_o_x_14[10];
  assign ofm_x_14_9 = uSystolicPE_388_io_ofm_d;
  assign randW_x_9_15 = uSystolicPE_388_io_randW_d;
  assign uSystolicPE_389_io_mac_done = mac_done_x_9[15];
  assign uSystolicPE_389_io_enable_i = enable_i_x_9[15];
  assign uSystolicPE_389_io_clear_i = clear_i_x_9[15];
  assign ifm_sign_x_9_16 = uSystolicPE_389_io_ifm_sign_d;
  assign ifm_dff_x_9_16 = uSystolicPE_389_io_ifm_dff_d;
  assign uSystolicPE_389_io_enable_w = enable_w_x_15[9];
  assign uSystolicPE_389_io_clear_w = clear_w_x_15[9];
  assign wght_sign_x_15_10 = uSystolicPE_389_io_wght_sign_d;
  assign wght_abs_x_15_10 = uSystolicPE_389_io_wght_abs_d;
  assign uSystolicPE_389_io_enable_o = enable_o_x_15[10];
  assign uSystolicPE_389_io_clear_o = clear_o_x_15[10];
  assign ofm_x_15_9 = uSystolicPE_389_io_ofm_d;
  assign randW_x_9_16 = uSystolicPE_389_io_randW_d;
  assign uSystolicPEBorder_26_io_mac_done = mac_done_x_10[0];
  assign uSystolicPEBorder_26_io_enable_i = enable_i_x_10[0];
  assign uSystolicPEBorder_26_io_clear_i = clear_i_x_10[0];
  assign ifm_sign_x_10_1 = uSystolicPEBorder_26_io_ifm_sign_d;
  assign ifm_dff_x_10_1 = uSystolicPEBorder_26_io_ifm_dff_d;
  assign uSystolicPEBorder_26_io_enable_w = enable_w_x_0[10];
  assign uSystolicPEBorder_26_io_clear_w = clear_w_x_0[10];
  assign wght_sign_x_0_11 = uSystolicPEBorder_26_io_wght_sign_d;
  assign wght_abs_x_0_11 = uSystolicPEBorder_26_io_wght_abs_d;
  assign uSystolicPEBorder_26_io_enable_o = enable_o_x_0[11];
  assign uSystolicPEBorder_26_io_clear_o = clear_o_x_0[11];
  assign ofm_x_0_10 = uSystolicPEBorder_26_io_ofm_d;
  assign randW_x_10_1 = uSystolicPEBorder_26_io_randW_d;
  assign uSystolicPE_390_io_mac_done = mac_done_x_10[1];
  assign uSystolicPE_390_io_enable_i = enable_i_x_10[1];
  assign uSystolicPE_390_io_clear_i = clear_i_x_10[1];
  assign ifm_sign_x_10_2 = uSystolicPE_390_io_ifm_sign_d;
  assign ifm_dff_x_10_2 = uSystolicPE_390_io_ifm_dff_d;
  assign uSystolicPE_390_io_enable_w = enable_w_x_1[10];
  assign uSystolicPE_390_io_clear_w = clear_w_x_1[10];
  assign wght_sign_x_1_11 = uSystolicPE_390_io_wght_sign_d;
  assign wght_abs_x_1_11 = uSystolicPE_390_io_wght_abs_d;
  assign uSystolicPE_390_io_enable_o = enable_o_x_1[11];
  assign uSystolicPE_390_io_clear_o = clear_o_x_1[11];
  assign ofm_x_1_10 = uSystolicPE_390_io_ofm_d;
  assign randW_x_10_2 = uSystolicPE_390_io_randW_d;
  assign uSystolicPE_391_io_mac_done = mac_done_x_10[2];
  assign uSystolicPE_391_io_enable_i = enable_i_x_10[2];
  assign uSystolicPE_391_io_clear_i = clear_i_x_10[2];
  assign ifm_sign_x_10_3 = uSystolicPE_391_io_ifm_sign_d;
  assign ifm_dff_x_10_3 = uSystolicPE_391_io_ifm_dff_d;
  assign uSystolicPE_391_io_enable_w = enable_w_x_2[10];
  assign uSystolicPE_391_io_clear_w = clear_w_x_2[10];
  assign wght_sign_x_2_11 = uSystolicPE_391_io_wght_sign_d;
  assign wght_abs_x_2_11 = uSystolicPE_391_io_wght_abs_d;
  assign uSystolicPE_391_io_enable_o = enable_o_x_2[11];
  assign uSystolicPE_391_io_clear_o = clear_o_x_2[11];
  assign ofm_x_2_10 = uSystolicPE_391_io_ofm_d;
  assign randW_x_10_3 = uSystolicPE_391_io_randW_d;
  assign uSystolicPE_392_io_mac_done = mac_done_x_10[3];
  assign uSystolicPE_392_io_enable_i = enable_i_x_10[3];
  assign uSystolicPE_392_io_clear_i = clear_i_x_10[3];
  assign ifm_sign_x_10_4 = uSystolicPE_392_io_ifm_sign_d;
  assign ifm_dff_x_10_4 = uSystolicPE_392_io_ifm_dff_d;
  assign uSystolicPE_392_io_enable_w = enable_w_x_3[10];
  assign uSystolicPE_392_io_clear_w = clear_w_x_3[10];
  assign wght_sign_x_3_11 = uSystolicPE_392_io_wght_sign_d;
  assign wght_abs_x_3_11 = uSystolicPE_392_io_wght_abs_d;
  assign uSystolicPE_392_io_enable_o = enable_o_x_3[11];
  assign uSystolicPE_392_io_clear_o = clear_o_x_3[11];
  assign ofm_x_3_10 = uSystolicPE_392_io_ofm_d;
  assign randW_x_10_4 = uSystolicPE_392_io_randW_d;
  assign uSystolicPE_393_io_mac_done = mac_done_x_10[4];
  assign uSystolicPE_393_io_enable_i = enable_i_x_10[4];
  assign uSystolicPE_393_io_clear_i = clear_i_x_10[4];
  assign ifm_sign_x_10_5 = uSystolicPE_393_io_ifm_sign_d;
  assign ifm_dff_x_10_5 = uSystolicPE_393_io_ifm_dff_d;
  assign uSystolicPE_393_io_enable_w = enable_w_x_4[10];
  assign uSystolicPE_393_io_clear_w = clear_w_x_4[10];
  assign wght_sign_x_4_11 = uSystolicPE_393_io_wght_sign_d;
  assign wght_abs_x_4_11 = uSystolicPE_393_io_wght_abs_d;
  assign uSystolicPE_393_io_enable_o = enable_o_x_4[11];
  assign uSystolicPE_393_io_clear_o = clear_o_x_4[11];
  assign ofm_x_4_10 = uSystolicPE_393_io_ofm_d;
  assign randW_x_10_5 = uSystolicPE_393_io_randW_d;
  assign uSystolicPE_394_io_mac_done = mac_done_x_10[5];
  assign uSystolicPE_394_io_enable_i = enable_i_x_10[5];
  assign uSystolicPE_394_io_clear_i = clear_i_x_10[5];
  assign ifm_sign_x_10_6 = uSystolicPE_394_io_ifm_sign_d;
  assign ifm_dff_x_10_6 = uSystolicPE_394_io_ifm_dff_d;
  assign uSystolicPE_394_io_enable_w = enable_w_x_5[10];
  assign uSystolicPE_394_io_clear_w = clear_w_x_5[10];
  assign wght_sign_x_5_11 = uSystolicPE_394_io_wght_sign_d;
  assign wght_abs_x_5_11 = uSystolicPE_394_io_wght_abs_d;
  assign uSystolicPE_394_io_enable_o = enable_o_x_5[11];
  assign uSystolicPE_394_io_clear_o = clear_o_x_5[11];
  assign ofm_x_5_10 = uSystolicPE_394_io_ofm_d;
  assign randW_x_10_6 = uSystolicPE_394_io_randW_d;
  assign uSystolicPE_395_io_mac_done = mac_done_x_10[6];
  assign uSystolicPE_395_io_enable_i = enable_i_x_10[6];
  assign uSystolicPE_395_io_clear_i = clear_i_x_10[6];
  assign ifm_sign_x_10_7 = uSystolicPE_395_io_ifm_sign_d;
  assign ifm_dff_x_10_7 = uSystolicPE_395_io_ifm_dff_d;
  assign uSystolicPE_395_io_enable_w = enable_w_x_6[10];
  assign uSystolicPE_395_io_clear_w = clear_w_x_6[10];
  assign wght_sign_x_6_11 = uSystolicPE_395_io_wght_sign_d;
  assign wght_abs_x_6_11 = uSystolicPE_395_io_wght_abs_d;
  assign uSystolicPE_395_io_enable_o = enable_o_x_6[11];
  assign uSystolicPE_395_io_clear_o = clear_o_x_6[11];
  assign ofm_x_6_10 = uSystolicPE_395_io_ofm_d;
  assign randW_x_10_7 = uSystolicPE_395_io_randW_d;
  assign uSystolicPE_396_io_mac_done = mac_done_x_10[7];
  assign uSystolicPE_396_io_enable_i = enable_i_x_10[7];
  assign uSystolicPE_396_io_clear_i = clear_i_x_10[7];
  assign ifm_sign_x_10_8 = uSystolicPE_396_io_ifm_sign_d;
  assign ifm_dff_x_10_8 = uSystolicPE_396_io_ifm_dff_d;
  assign uSystolicPE_396_io_enable_w = enable_w_x_7[10];
  assign uSystolicPE_396_io_clear_w = clear_w_x_7[10];
  assign wght_sign_x_7_11 = uSystolicPE_396_io_wght_sign_d;
  assign wght_abs_x_7_11 = uSystolicPE_396_io_wght_abs_d;
  assign uSystolicPE_396_io_enable_o = enable_o_x_7[11];
  assign uSystolicPE_396_io_clear_o = clear_o_x_7[11];
  assign ofm_x_7_10 = uSystolicPE_396_io_ofm_d;
  assign randW_x_10_8 = uSystolicPE_396_io_randW_d;
  assign uSystolicPE_397_io_mac_done = mac_done_x_10[8];
  assign uSystolicPE_397_io_enable_i = enable_i_x_10[8];
  assign uSystolicPE_397_io_clear_i = clear_i_x_10[8];
  assign ifm_sign_x_10_9 = uSystolicPE_397_io_ifm_sign_d;
  assign ifm_dff_x_10_9 = uSystolicPE_397_io_ifm_dff_d;
  assign uSystolicPE_397_io_enable_w = enable_w_x_8[10];
  assign uSystolicPE_397_io_clear_w = clear_w_x_8[10];
  assign wght_sign_x_8_11 = uSystolicPE_397_io_wght_sign_d;
  assign wght_abs_x_8_11 = uSystolicPE_397_io_wght_abs_d;
  assign uSystolicPE_397_io_enable_o = enable_o_x_8[11];
  assign uSystolicPE_397_io_clear_o = clear_o_x_8[11];
  assign ofm_x_8_10 = uSystolicPE_397_io_ofm_d;
  assign randW_x_10_9 = uSystolicPE_397_io_randW_d;
  assign uSystolicPE_398_io_mac_done = mac_done_x_10[9];
  assign uSystolicPE_398_io_enable_i = enable_i_x_10[9];
  assign uSystolicPE_398_io_clear_i = clear_i_x_10[9];
  assign ifm_sign_x_10_10 = uSystolicPE_398_io_ifm_sign_d;
  assign ifm_dff_x_10_10 = uSystolicPE_398_io_ifm_dff_d;
  assign uSystolicPE_398_io_enable_w = enable_w_x_9[10];
  assign uSystolicPE_398_io_clear_w = clear_w_x_9[10];
  assign wght_sign_x_9_11 = uSystolicPE_398_io_wght_sign_d;
  assign wght_abs_x_9_11 = uSystolicPE_398_io_wght_abs_d;
  assign uSystolicPE_398_io_enable_o = enable_o_x_9[11];
  assign uSystolicPE_398_io_clear_o = clear_o_x_9[11];
  assign ofm_x_9_10 = uSystolicPE_398_io_ofm_d;
  assign randW_x_10_10 = uSystolicPE_398_io_randW_d;
  assign uSystolicPE_399_io_mac_done = mac_done_x_10[10];
  assign uSystolicPE_399_io_enable_i = enable_i_x_10[10];
  assign uSystolicPE_399_io_clear_i = clear_i_x_10[10];
  assign ifm_sign_x_10_11 = uSystolicPE_399_io_ifm_sign_d;
  assign ifm_dff_x_10_11 = uSystolicPE_399_io_ifm_dff_d;
  assign uSystolicPE_399_io_enable_w = enable_w_x_10[10];
  assign uSystolicPE_399_io_clear_w = clear_w_x_10[10];
  assign wght_sign_x_10_11 = uSystolicPE_399_io_wght_sign_d;
  assign wght_abs_x_10_11 = uSystolicPE_399_io_wght_abs_d;
  assign uSystolicPE_399_io_enable_o = enable_o_x_10[11];
  assign uSystolicPE_399_io_clear_o = clear_o_x_10[11];
  assign ofm_x_10_10 = uSystolicPE_399_io_ofm_d;
  assign randW_x_10_11 = uSystolicPE_399_io_randW_d;
  assign uSystolicPE_400_io_mac_done = mac_done_x_10[11];
  assign uSystolicPE_400_io_enable_i = enable_i_x_10[11];
  assign uSystolicPE_400_io_clear_i = clear_i_x_10[11];
  assign ifm_sign_x_10_12 = uSystolicPE_400_io_ifm_sign_d;
  assign ifm_dff_x_10_12 = uSystolicPE_400_io_ifm_dff_d;
  assign uSystolicPE_400_io_enable_w = enable_w_x_11[10];
  assign uSystolicPE_400_io_clear_w = clear_w_x_11[10];
  assign wght_sign_x_11_11 = uSystolicPE_400_io_wght_sign_d;
  assign wght_abs_x_11_11 = uSystolicPE_400_io_wght_abs_d;
  assign uSystolicPE_400_io_enable_o = enable_o_x_11[11];
  assign uSystolicPE_400_io_clear_o = clear_o_x_11[11];
  assign ofm_x_11_10 = uSystolicPE_400_io_ofm_d;
  assign randW_x_10_12 = uSystolicPE_400_io_randW_d;
  assign uSystolicPE_401_io_mac_done = mac_done_x_10[12];
  assign uSystolicPE_401_io_enable_i = enable_i_x_10[12];
  assign uSystolicPE_401_io_clear_i = clear_i_x_10[12];
  assign ifm_sign_x_10_13 = uSystolicPE_401_io_ifm_sign_d;
  assign ifm_dff_x_10_13 = uSystolicPE_401_io_ifm_dff_d;
  assign uSystolicPE_401_io_enable_w = enable_w_x_12[10];
  assign uSystolicPE_401_io_clear_w = clear_w_x_12[10];
  assign wght_sign_x_12_11 = uSystolicPE_401_io_wght_sign_d;
  assign wght_abs_x_12_11 = uSystolicPE_401_io_wght_abs_d;
  assign uSystolicPE_401_io_enable_o = enable_o_x_12[11];
  assign uSystolicPE_401_io_clear_o = clear_o_x_12[11];
  assign ofm_x_12_10 = uSystolicPE_401_io_ofm_d;
  assign randW_x_10_13 = uSystolicPE_401_io_randW_d;
  assign uSystolicPE_402_io_mac_done = mac_done_x_10[13];
  assign uSystolicPE_402_io_enable_i = enable_i_x_10[13];
  assign uSystolicPE_402_io_clear_i = clear_i_x_10[13];
  assign ifm_sign_x_10_14 = uSystolicPE_402_io_ifm_sign_d;
  assign ifm_dff_x_10_14 = uSystolicPE_402_io_ifm_dff_d;
  assign uSystolicPE_402_io_enable_w = enable_w_x_13[10];
  assign uSystolicPE_402_io_clear_w = clear_w_x_13[10];
  assign wght_sign_x_13_11 = uSystolicPE_402_io_wght_sign_d;
  assign wght_abs_x_13_11 = uSystolicPE_402_io_wght_abs_d;
  assign uSystolicPE_402_io_enable_o = enable_o_x_13[11];
  assign uSystolicPE_402_io_clear_o = clear_o_x_13[11];
  assign ofm_x_13_10 = uSystolicPE_402_io_ofm_d;
  assign randW_x_10_14 = uSystolicPE_402_io_randW_d;
  assign uSystolicPE_403_io_mac_done = mac_done_x_10[14];
  assign uSystolicPE_403_io_enable_i = enable_i_x_10[14];
  assign uSystolicPE_403_io_clear_i = clear_i_x_10[14];
  assign ifm_sign_x_10_15 = uSystolicPE_403_io_ifm_sign_d;
  assign ifm_dff_x_10_15 = uSystolicPE_403_io_ifm_dff_d;
  assign uSystolicPE_403_io_enable_w = enable_w_x_14[10];
  assign uSystolicPE_403_io_clear_w = clear_w_x_14[10];
  assign wght_sign_x_14_11 = uSystolicPE_403_io_wght_sign_d;
  assign wght_abs_x_14_11 = uSystolicPE_403_io_wght_abs_d;
  assign uSystolicPE_403_io_enable_o = enable_o_x_14[11];
  assign uSystolicPE_403_io_clear_o = clear_o_x_14[11];
  assign ofm_x_14_10 = uSystolicPE_403_io_ofm_d;
  assign randW_x_10_15 = uSystolicPE_403_io_randW_d;
  assign uSystolicPE_404_io_mac_done = mac_done_x_10[15];
  assign uSystolicPE_404_io_enable_i = enable_i_x_10[15];
  assign uSystolicPE_404_io_clear_i = clear_i_x_10[15];
  assign ifm_sign_x_10_16 = uSystolicPE_404_io_ifm_sign_d;
  assign ifm_dff_x_10_16 = uSystolicPE_404_io_ifm_dff_d;
  assign uSystolicPE_404_io_enable_w = enable_w_x_15[10];
  assign uSystolicPE_404_io_clear_w = clear_w_x_15[10];
  assign wght_sign_x_15_11 = uSystolicPE_404_io_wght_sign_d;
  assign wght_abs_x_15_11 = uSystolicPE_404_io_wght_abs_d;
  assign uSystolicPE_404_io_enable_o = enable_o_x_15[11];
  assign uSystolicPE_404_io_clear_o = clear_o_x_15[11];
  assign ofm_x_15_10 = uSystolicPE_404_io_ofm_d;
  assign randW_x_10_16 = uSystolicPE_404_io_randW_d;
  assign uSystolicPEBorder_27_io_mac_done = mac_done_x_11[0];
  assign uSystolicPEBorder_27_io_enable_i = enable_i_x_11[0];
  assign uSystolicPEBorder_27_io_clear_i = clear_i_x_11[0];
  assign ifm_sign_x_11_1 = uSystolicPEBorder_27_io_ifm_sign_d;
  assign ifm_dff_x_11_1 = uSystolicPEBorder_27_io_ifm_dff_d;
  assign uSystolicPEBorder_27_io_enable_w = enable_w_x_0[11];
  assign uSystolicPEBorder_27_io_clear_w = clear_w_x_0[11];
  assign wght_sign_x_0_12 = uSystolicPEBorder_27_io_wght_sign_d;
  assign wght_abs_x_0_12 = uSystolicPEBorder_27_io_wght_abs_d;
  assign uSystolicPEBorder_27_io_enable_o = enable_o_x_0[12];
  assign uSystolicPEBorder_27_io_clear_o = clear_o_x_0[12];
  assign ofm_x_0_11 = uSystolicPEBorder_27_io_ofm_d;
  assign randW_x_11_1 = uSystolicPEBorder_27_io_randW_d;
  assign uSystolicPE_405_io_mac_done = mac_done_x_11[1];
  assign uSystolicPE_405_io_enable_i = enable_i_x_11[1];
  assign uSystolicPE_405_io_clear_i = clear_i_x_11[1];
  assign ifm_sign_x_11_2 = uSystolicPE_405_io_ifm_sign_d;
  assign ifm_dff_x_11_2 = uSystolicPE_405_io_ifm_dff_d;
  assign uSystolicPE_405_io_enable_w = enable_w_x_1[11];
  assign uSystolicPE_405_io_clear_w = clear_w_x_1[11];
  assign wght_sign_x_1_12 = uSystolicPE_405_io_wght_sign_d;
  assign wght_abs_x_1_12 = uSystolicPE_405_io_wght_abs_d;
  assign uSystolicPE_405_io_enable_o = enable_o_x_1[12];
  assign uSystolicPE_405_io_clear_o = clear_o_x_1[12];
  assign ofm_x_1_11 = uSystolicPE_405_io_ofm_d;
  assign randW_x_11_2 = uSystolicPE_405_io_randW_d;
  assign uSystolicPE_406_io_mac_done = mac_done_x_11[2];
  assign uSystolicPE_406_io_enable_i = enable_i_x_11[2];
  assign uSystolicPE_406_io_clear_i = clear_i_x_11[2];
  assign ifm_sign_x_11_3 = uSystolicPE_406_io_ifm_sign_d;
  assign ifm_dff_x_11_3 = uSystolicPE_406_io_ifm_dff_d;
  assign uSystolicPE_406_io_enable_w = enable_w_x_2[11];
  assign uSystolicPE_406_io_clear_w = clear_w_x_2[11];
  assign wght_sign_x_2_12 = uSystolicPE_406_io_wght_sign_d;
  assign wght_abs_x_2_12 = uSystolicPE_406_io_wght_abs_d;
  assign uSystolicPE_406_io_enable_o = enable_o_x_2[12];
  assign uSystolicPE_406_io_clear_o = clear_o_x_2[12];
  assign ofm_x_2_11 = uSystolicPE_406_io_ofm_d;
  assign randW_x_11_3 = uSystolicPE_406_io_randW_d;
  assign uSystolicPE_407_io_mac_done = mac_done_x_11[3];
  assign uSystolicPE_407_io_enable_i = enable_i_x_11[3];
  assign uSystolicPE_407_io_clear_i = clear_i_x_11[3];
  assign ifm_sign_x_11_4 = uSystolicPE_407_io_ifm_sign_d;
  assign ifm_dff_x_11_4 = uSystolicPE_407_io_ifm_dff_d;
  assign uSystolicPE_407_io_enable_w = enable_w_x_3[11];
  assign uSystolicPE_407_io_clear_w = clear_w_x_3[11];
  assign wght_sign_x_3_12 = uSystolicPE_407_io_wght_sign_d;
  assign wght_abs_x_3_12 = uSystolicPE_407_io_wght_abs_d;
  assign uSystolicPE_407_io_enable_o = enable_o_x_3[12];
  assign uSystolicPE_407_io_clear_o = clear_o_x_3[12];
  assign ofm_x_3_11 = uSystolicPE_407_io_ofm_d;
  assign randW_x_11_4 = uSystolicPE_407_io_randW_d;
  assign uSystolicPE_408_io_mac_done = mac_done_x_11[4];
  assign uSystolicPE_408_io_enable_i = enable_i_x_11[4];
  assign uSystolicPE_408_io_clear_i = clear_i_x_11[4];
  assign ifm_sign_x_11_5 = uSystolicPE_408_io_ifm_sign_d;
  assign ifm_dff_x_11_5 = uSystolicPE_408_io_ifm_dff_d;
  assign uSystolicPE_408_io_enable_w = enable_w_x_4[11];
  assign uSystolicPE_408_io_clear_w = clear_w_x_4[11];
  assign wght_sign_x_4_12 = uSystolicPE_408_io_wght_sign_d;
  assign wght_abs_x_4_12 = uSystolicPE_408_io_wght_abs_d;
  assign uSystolicPE_408_io_enable_o = enable_o_x_4[12];
  assign uSystolicPE_408_io_clear_o = clear_o_x_4[12];
  assign ofm_x_4_11 = uSystolicPE_408_io_ofm_d;
  assign randW_x_11_5 = uSystolicPE_408_io_randW_d;
  assign uSystolicPE_409_io_mac_done = mac_done_x_11[5];
  assign uSystolicPE_409_io_enable_i = enable_i_x_11[5];
  assign uSystolicPE_409_io_clear_i = clear_i_x_11[5];
  assign ifm_sign_x_11_6 = uSystolicPE_409_io_ifm_sign_d;
  assign ifm_dff_x_11_6 = uSystolicPE_409_io_ifm_dff_d;
  assign uSystolicPE_409_io_enable_w = enable_w_x_5[11];
  assign uSystolicPE_409_io_clear_w = clear_w_x_5[11];
  assign wght_sign_x_5_12 = uSystolicPE_409_io_wght_sign_d;
  assign wght_abs_x_5_12 = uSystolicPE_409_io_wght_abs_d;
  assign uSystolicPE_409_io_enable_o = enable_o_x_5[12];
  assign uSystolicPE_409_io_clear_o = clear_o_x_5[12];
  assign ofm_x_5_11 = uSystolicPE_409_io_ofm_d;
  assign randW_x_11_6 = uSystolicPE_409_io_randW_d;
  assign uSystolicPE_410_io_mac_done = mac_done_x_11[6];
  assign uSystolicPE_410_io_enable_i = enable_i_x_11[6];
  assign uSystolicPE_410_io_clear_i = clear_i_x_11[6];
  assign ifm_sign_x_11_7 = uSystolicPE_410_io_ifm_sign_d;
  assign ifm_dff_x_11_7 = uSystolicPE_410_io_ifm_dff_d;
  assign uSystolicPE_410_io_enable_w = enable_w_x_6[11];
  assign uSystolicPE_410_io_clear_w = clear_w_x_6[11];
  assign wght_sign_x_6_12 = uSystolicPE_410_io_wght_sign_d;
  assign wght_abs_x_6_12 = uSystolicPE_410_io_wght_abs_d;
  assign uSystolicPE_410_io_enable_o = enable_o_x_6[12];
  assign uSystolicPE_410_io_clear_o = clear_o_x_6[12];
  assign ofm_x_6_11 = uSystolicPE_410_io_ofm_d;
  assign randW_x_11_7 = uSystolicPE_410_io_randW_d;
  assign uSystolicPE_411_io_mac_done = mac_done_x_11[7];
  assign uSystolicPE_411_io_enable_i = enable_i_x_11[7];
  assign uSystolicPE_411_io_clear_i = clear_i_x_11[7];
  assign ifm_sign_x_11_8 = uSystolicPE_411_io_ifm_sign_d;
  assign ifm_dff_x_11_8 = uSystolicPE_411_io_ifm_dff_d;
  assign uSystolicPE_411_io_enable_w = enable_w_x_7[11];
  assign uSystolicPE_411_io_clear_w = clear_w_x_7[11];
  assign wght_sign_x_7_12 = uSystolicPE_411_io_wght_sign_d;
  assign wght_abs_x_7_12 = uSystolicPE_411_io_wght_abs_d;
  assign uSystolicPE_411_io_enable_o = enable_o_x_7[12];
  assign uSystolicPE_411_io_clear_o = clear_o_x_7[12];
  assign ofm_x_7_11 = uSystolicPE_411_io_ofm_d;
  assign randW_x_11_8 = uSystolicPE_411_io_randW_d;
  assign uSystolicPE_412_io_mac_done = mac_done_x_11[8];
  assign uSystolicPE_412_io_enable_i = enable_i_x_11[8];
  assign uSystolicPE_412_io_clear_i = clear_i_x_11[8];
  assign ifm_sign_x_11_9 = uSystolicPE_412_io_ifm_sign_d;
  assign ifm_dff_x_11_9 = uSystolicPE_412_io_ifm_dff_d;
  assign uSystolicPE_412_io_enable_w = enable_w_x_8[11];
  assign uSystolicPE_412_io_clear_w = clear_w_x_8[11];
  assign wght_sign_x_8_12 = uSystolicPE_412_io_wght_sign_d;
  assign wght_abs_x_8_12 = uSystolicPE_412_io_wght_abs_d;
  assign uSystolicPE_412_io_enable_o = enable_o_x_8[12];
  assign uSystolicPE_412_io_clear_o = clear_o_x_8[12];
  assign ofm_x_8_11 = uSystolicPE_412_io_ofm_d;
  assign randW_x_11_9 = uSystolicPE_412_io_randW_d;
  assign uSystolicPE_413_io_mac_done = mac_done_x_11[9];
  assign uSystolicPE_413_io_enable_i = enable_i_x_11[9];
  assign uSystolicPE_413_io_clear_i = clear_i_x_11[9];
  assign ifm_sign_x_11_10 = uSystolicPE_413_io_ifm_sign_d;
  assign ifm_dff_x_11_10 = uSystolicPE_413_io_ifm_dff_d;
  assign uSystolicPE_413_io_enable_w = enable_w_x_9[11];
  assign uSystolicPE_413_io_clear_w = clear_w_x_9[11];
  assign wght_sign_x_9_12 = uSystolicPE_413_io_wght_sign_d;
  assign wght_abs_x_9_12 = uSystolicPE_413_io_wght_abs_d;
  assign uSystolicPE_413_io_enable_o = enable_o_x_9[12];
  assign uSystolicPE_413_io_clear_o = clear_o_x_9[12];
  assign ofm_x_9_11 = uSystolicPE_413_io_ofm_d;
  assign randW_x_11_10 = uSystolicPE_413_io_randW_d;
  assign uSystolicPE_414_io_mac_done = mac_done_x_11[10];
  assign uSystolicPE_414_io_enable_i = enable_i_x_11[10];
  assign uSystolicPE_414_io_clear_i = clear_i_x_11[10];
  assign ifm_sign_x_11_11 = uSystolicPE_414_io_ifm_sign_d;
  assign ifm_dff_x_11_11 = uSystolicPE_414_io_ifm_dff_d;
  assign uSystolicPE_414_io_enable_w = enable_w_x_10[11];
  assign uSystolicPE_414_io_clear_w = clear_w_x_10[11];
  assign wght_sign_x_10_12 = uSystolicPE_414_io_wght_sign_d;
  assign wght_abs_x_10_12 = uSystolicPE_414_io_wght_abs_d;
  assign uSystolicPE_414_io_enable_o = enable_o_x_10[12];
  assign uSystolicPE_414_io_clear_o = clear_o_x_10[12];
  assign ofm_x_10_11 = uSystolicPE_414_io_ofm_d;
  assign randW_x_11_11 = uSystolicPE_414_io_randW_d;
  assign uSystolicPE_415_io_mac_done = mac_done_x_11[11];
  assign uSystolicPE_415_io_enable_i = enable_i_x_11[11];
  assign uSystolicPE_415_io_clear_i = clear_i_x_11[11];
  assign ifm_sign_x_11_12 = uSystolicPE_415_io_ifm_sign_d;
  assign ifm_dff_x_11_12 = uSystolicPE_415_io_ifm_dff_d;
  assign uSystolicPE_415_io_enable_w = enable_w_x_11[11];
  assign uSystolicPE_415_io_clear_w = clear_w_x_11[11];
  assign wght_sign_x_11_12 = uSystolicPE_415_io_wght_sign_d;
  assign wght_abs_x_11_12 = uSystolicPE_415_io_wght_abs_d;
  assign uSystolicPE_415_io_enable_o = enable_o_x_11[12];
  assign uSystolicPE_415_io_clear_o = clear_o_x_11[12];
  assign ofm_x_11_11 = uSystolicPE_415_io_ofm_d;
  assign randW_x_11_12 = uSystolicPE_415_io_randW_d;
  assign uSystolicPE_416_io_mac_done = mac_done_x_11[12];
  assign uSystolicPE_416_io_enable_i = enable_i_x_11[12];
  assign uSystolicPE_416_io_clear_i = clear_i_x_11[12];
  assign ifm_sign_x_11_13 = uSystolicPE_416_io_ifm_sign_d;
  assign ifm_dff_x_11_13 = uSystolicPE_416_io_ifm_dff_d;
  assign uSystolicPE_416_io_enable_w = enable_w_x_12[11];
  assign uSystolicPE_416_io_clear_w = clear_w_x_12[11];
  assign wght_sign_x_12_12 = uSystolicPE_416_io_wght_sign_d;
  assign wght_abs_x_12_12 = uSystolicPE_416_io_wght_abs_d;
  assign uSystolicPE_416_io_enable_o = enable_o_x_12[12];
  assign uSystolicPE_416_io_clear_o = clear_o_x_12[12];
  assign ofm_x_12_11 = uSystolicPE_416_io_ofm_d;
  assign randW_x_11_13 = uSystolicPE_416_io_randW_d;
  assign uSystolicPE_417_io_mac_done = mac_done_x_11[13];
  assign uSystolicPE_417_io_enable_i = enable_i_x_11[13];
  assign uSystolicPE_417_io_clear_i = clear_i_x_11[13];
  assign ifm_sign_x_11_14 = uSystolicPE_417_io_ifm_sign_d;
  assign ifm_dff_x_11_14 = uSystolicPE_417_io_ifm_dff_d;
  assign uSystolicPE_417_io_enable_w = enable_w_x_13[11];
  assign uSystolicPE_417_io_clear_w = clear_w_x_13[11];
  assign wght_sign_x_13_12 = uSystolicPE_417_io_wght_sign_d;
  assign wght_abs_x_13_12 = uSystolicPE_417_io_wght_abs_d;
  assign uSystolicPE_417_io_enable_o = enable_o_x_13[12];
  assign uSystolicPE_417_io_clear_o = clear_o_x_13[12];
  assign ofm_x_13_11 = uSystolicPE_417_io_ofm_d;
  assign randW_x_11_14 = uSystolicPE_417_io_randW_d;
  assign uSystolicPE_418_io_mac_done = mac_done_x_11[14];
  assign uSystolicPE_418_io_enable_i = enable_i_x_11[14];
  assign uSystolicPE_418_io_clear_i = clear_i_x_11[14];
  assign ifm_sign_x_11_15 = uSystolicPE_418_io_ifm_sign_d;
  assign ifm_dff_x_11_15 = uSystolicPE_418_io_ifm_dff_d;
  assign uSystolicPE_418_io_enable_w = enable_w_x_14[11];
  assign uSystolicPE_418_io_clear_w = clear_w_x_14[11];
  assign wght_sign_x_14_12 = uSystolicPE_418_io_wght_sign_d;
  assign wght_abs_x_14_12 = uSystolicPE_418_io_wght_abs_d;
  assign uSystolicPE_418_io_enable_o = enable_o_x_14[12];
  assign uSystolicPE_418_io_clear_o = clear_o_x_14[12];
  assign ofm_x_14_11 = uSystolicPE_418_io_ofm_d;
  assign randW_x_11_15 = uSystolicPE_418_io_randW_d;
  assign uSystolicPE_419_io_mac_done = mac_done_x_11[15];
  assign uSystolicPE_419_io_enable_i = enable_i_x_11[15];
  assign uSystolicPE_419_io_clear_i = clear_i_x_11[15];
  assign ifm_sign_x_11_16 = uSystolicPE_419_io_ifm_sign_d;
  assign ifm_dff_x_11_16 = uSystolicPE_419_io_ifm_dff_d;
  assign uSystolicPE_419_io_enable_w = enable_w_x_15[11];
  assign uSystolicPE_419_io_clear_w = clear_w_x_15[11];
  assign wght_sign_x_15_12 = uSystolicPE_419_io_wght_sign_d;
  assign wght_abs_x_15_12 = uSystolicPE_419_io_wght_abs_d;
  assign uSystolicPE_419_io_enable_o = enable_o_x_15[12];
  assign uSystolicPE_419_io_clear_o = clear_o_x_15[12];
  assign ofm_x_15_11 = uSystolicPE_419_io_ofm_d;
  assign randW_x_11_16 = uSystolicPE_419_io_randW_d;
  assign uSystolicPEBorder_28_io_mac_done = mac_done_x_12[0];
  assign uSystolicPEBorder_28_io_enable_i = enable_i_x_12[0];
  assign uSystolicPEBorder_28_io_clear_i = clear_i_x_12[0];
  assign ifm_sign_x_12_1 = uSystolicPEBorder_28_io_ifm_sign_d;
  assign ifm_dff_x_12_1 = uSystolicPEBorder_28_io_ifm_dff_d;
  assign uSystolicPEBorder_28_io_enable_w = enable_w_x_0[12];
  assign uSystolicPEBorder_28_io_clear_w = clear_w_x_0[12];
  assign wght_sign_x_0_13 = uSystolicPEBorder_28_io_wght_sign_d;
  assign wght_abs_x_0_13 = uSystolicPEBorder_28_io_wght_abs_d;
  assign uSystolicPEBorder_28_io_enable_o = enable_o_x_0[13];
  assign uSystolicPEBorder_28_io_clear_o = clear_o_x_0[13];
  assign ofm_x_0_12 = uSystolicPEBorder_28_io_ofm_d;
  assign randW_x_12_1 = uSystolicPEBorder_28_io_randW_d;
  assign uSystolicPE_420_io_mac_done = mac_done_x_12[1];
  assign uSystolicPE_420_io_enable_i = enable_i_x_12[1];
  assign uSystolicPE_420_io_clear_i = clear_i_x_12[1];
  assign ifm_sign_x_12_2 = uSystolicPE_420_io_ifm_sign_d;
  assign ifm_dff_x_12_2 = uSystolicPE_420_io_ifm_dff_d;
  assign uSystolicPE_420_io_enable_w = enable_w_x_1[12];
  assign uSystolicPE_420_io_clear_w = clear_w_x_1[12];
  assign wght_sign_x_1_13 = uSystolicPE_420_io_wght_sign_d;
  assign wght_abs_x_1_13 = uSystolicPE_420_io_wght_abs_d;
  assign uSystolicPE_420_io_enable_o = enable_o_x_1[13];
  assign uSystolicPE_420_io_clear_o = clear_o_x_1[13];
  assign ofm_x_1_12 = uSystolicPE_420_io_ofm_d;
  assign randW_x_12_2 = uSystolicPE_420_io_randW_d;
  assign uSystolicPE_421_io_mac_done = mac_done_x_12[2];
  assign uSystolicPE_421_io_enable_i = enable_i_x_12[2];
  assign uSystolicPE_421_io_clear_i = clear_i_x_12[2];
  assign ifm_sign_x_12_3 = uSystolicPE_421_io_ifm_sign_d;
  assign ifm_dff_x_12_3 = uSystolicPE_421_io_ifm_dff_d;
  assign uSystolicPE_421_io_enable_w = enable_w_x_2[12];
  assign uSystolicPE_421_io_clear_w = clear_w_x_2[12];
  assign wght_sign_x_2_13 = uSystolicPE_421_io_wght_sign_d;
  assign wght_abs_x_2_13 = uSystolicPE_421_io_wght_abs_d;
  assign uSystolicPE_421_io_enable_o = enable_o_x_2[13];
  assign uSystolicPE_421_io_clear_o = clear_o_x_2[13];
  assign ofm_x_2_12 = uSystolicPE_421_io_ofm_d;
  assign randW_x_12_3 = uSystolicPE_421_io_randW_d;
  assign uSystolicPE_422_io_mac_done = mac_done_x_12[3];
  assign uSystolicPE_422_io_enable_i = enable_i_x_12[3];
  assign uSystolicPE_422_io_clear_i = clear_i_x_12[3];
  assign ifm_sign_x_12_4 = uSystolicPE_422_io_ifm_sign_d;
  assign ifm_dff_x_12_4 = uSystolicPE_422_io_ifm_dff_d;
  assign uSystolicPE_422_io_enable_w = enable_w_x_3[12];
  assign uSystolicPE_422_io_clear_w = clear_w_x_3[12];
  assign wght_sign_x_3_13 = uSystolicPE_422_io_wght_sign_d;
  assign wght_abs_x_3_13 = uSystolicPE_422_io_wght_abs_d;
  assign uSystolicPE_422_io_enable_o = enable_o_x_3[13];
  assign uSystolicPE_422_io_clear_o = clear_o_x_3[13];
  assign ofm_x_3_12 = uSystolicPE_422_io_ofm_d;
  assign randW_x_12_4 = uSystolicPE_422_io_randW_d;
  assign uSystolicPE_423_io_mac_done = mac_done_x_12[4];
  assign uSystolicPE_423_io_enable_i = enable_i_x_12[4];
  assign uSystolicPE_423_io_clear_i = clear_i_x_12[4];
  assign ifm_sign_x_12_5 = uSystolicPE_423_io_ifm_sign_d;
  assign ifm_dff_x_12_5 = uSystolicPE_423_io_ifm_dff_d;
  assign uSystolicPE_423_io_enable_w = enable_w_x_4[12];
  assign uSystolicPE_423_io_clear_w = clear_w_x_4[12];
  assign wght_sign_x_4_13 = uSystolicPE_423_io_wght_sign_d;
  assign wght_abs_x_4_13 = uSystolicPE_423_io_wght_abs_d;
  assign uSystolicPE_423_io_enable_o = enable_o_x_4[13];
  assign uSystolicPE_423_io_clear_o = clear_o_x_4[13];
  assign ofm_x_4_12 = uSystolicPE_423_io_ofm_d;
  assign randW_x_12_5 = uSystolicPE_423_io_randW_d;
  assign uSystolicPE_424_io_mac_done = mac_done_x_12[5];
  assign uSystolicPE_424_io_enable_i = enable_i_x_12[5];
  assign uSystolicPE_424_io_clear_i = clear_i_x_12[5];
  assign ifm_sign_x_12_6 = uSystolicPE_424_io_ifm_sign_d;
  assign ifm_dff_x_12_6 = uSystolicPE_424_io_ifm_dff_d;
  assign uSystolicPE_424_io_enable_w = enable_w_x_5[12];
  assign uSystolicPE_424_io_clear_w = clear_w_x_5[12];
  assign wght_sign_x_5_13 = uSystolicPE_424_io_wght_sign_d;
  assign wght_abs_x_5_13 = uSystolicPE_424_io_wght_abs_d;
  assign uSystolicPE_424_io_enable_o = enable_o_x_5[13];
  assign uSystolicPE_424_io_clear_o = clear_o_x_5[13];
  assign ofm_x_5_12 = uSystolicPE_424_io_ofm_d;
  assign randW_x_12_6 = uSystolicPE_424_io_randW_d;
  assign uSystolicPE_425_io_mac_done = mac_done_x_12[6];
  assign uSystolicPE_425_io_enable_i = enable_i_x_12[6];
  assign uSystolicPE_425_io_clear_i = clear_i_x_12[6];
  assign ifm_sign_x_12_7 = uSystolicPE_425_io_ifm_sign_d;
  assign ifm_dff_x_12_7 = uSystolicPE_425_io_ifm_dff_d;
  assign uSystolicPE_425_io_enable_w = enable_w_x_6[12];
  assign uSystolicPE_425_io_clear_w = clear_w_x_6[12];
  assign wght_sign_x_6_13 = uSystolicPE_425_io_wght_sign_d;
  assign wght_abs_x_6_13 = uSystolicPE_425_io_wght_abs_d;
  assign uSystolicPE_425_io_enable_o = enable_o_x_6[13];
  assign uSystolicPE_425_io_clear_o = clear_o_x_6[13];
  assign ofm_x_6_12 = uSystolicPE_425_io_ofm_d;
  assign randW_x_12_7 = uSystolicPE_425_io_randW_d;
  assign uSystolicPE_426_io_mac_done = mac_done_x_12[7];
  assign uSystolicPE_426_io_enable_i = enable_i_x_12[7];
  assign uSystolicPE_426_io_clear_i = clear_i_x_12[7];
  assign ifm_sign_x_12_8 = uSystolicPE_426_io_ifm_sign_d;
  assign ifm_dff_x_12_8 = uSystolicPE_426_io_ifm_dff_d;
  assign uSystolicPE_426_io_enable_w = enable_w_x_7[12];
  assign uSystolicPE_426_io_clear_w = clear_w_x_7[12];
  assign wght_sign_x_7_13 = uSystolicPE_426_io_wght_sign_d;
  assign wght_abs_x_7_13 = uSystolicPE_426_io_wght_abs_d;
  assign uSystolicPE_426_io_enable_o = enable_o_x_7[13];
  assign uSystolicPE_426_io_clear_o = clear_o_x_7[13];
  assign ofm_x_7_12 = uSystolicPE_426_io_ofm_d;
  assign randW_x_12_8 = uSystolicPE_426_io_randW_d;
  assign uSystolicPE_427_io_mac_done = mac_done_x_12[8];
  assign uSystolicPE_427_io_enable_i = enable_i_x_12[8];
  assign uSystolicPE_427_io_clear_i = clear_i_x_12[8];
  assign ifm_sign_x_12_9 = uSystolicPE_427_io_ifm_sign_d;
  assign ifm_dff_x_12_9 = uSystolicPE_427_io_ifm_dff_d;
  assign uSystolicPE_427_io_enable_w = enable_w_x_8[12];
  assign uSystolicPE_427_io_clear_w = clear_w_x_8[12];
  assign wght_sign_x_8_13 = uSystolicPE_427_io_wght_sign_d;
  assign wght_abs_x_8_13 = uSystolicPE_427_io_wght_abs_d;
  assign uSystolicPE_427_io_enable_o = enable_o_x_8[13];
  assign uSystolicPE_427_io_clear_o = clear_o_x_8[13];
  assign ofm_x_8_12 = uSystolicPE_427_io_ofm_d;
  assign randW_x_12_9 = uSystolicPE_427_io_randW_d;
  assign uSystolicPE_428_io_mac_done = mac_done_x_12[9];
  assign uSystolicPE_428_io_enable_i = enable_i_x_12[9];
  assign uSystolicPE_428_io_clear_i = clear_i_x_12[9];
  assign ifm_sign_x_12_10 = uSystolicPE_428_io_ifm_sign_d;
  assign ifm_dff_x_12_10 = uSystolicPE_428_io_ifm_dff_d;
  assign uSystolicPE_428_io_enable_w = enable_w_x_9[12];
  assign uSystolicPE_428_io_clear_w = clear_w_x_9[12];
  assign wght_sign_x_9_13 = uSystolicPE_428_io_wght_sign_d;
  assign wght_abs_x_9_13 = uSystolicPE_428_io_wght_abs_d;
  assign uSystolicPE_428_io_enable_o = enable_o_x_9[13];
  assign uSystolicPE_428_io_clear_o = clear_o_x_9[13];
  assign ofm_x_9_12 = uSystolicPE_428_io_ofm_d;
  assign randW_x_12_10 = uSystolicPE_428_io_randW_d;
  assign uSystolicPE_429_io_mac_done = mac_done_x_12[10];
  assign uSystolicPE_429_io_enable_i = enable_i_x_12[10];
  assign uSystolicPE_429_io_clear_i = clear_i_x_12[10];
  assign ifm_sign_x_12_11 = uSystolicPE_429_io_ifm_sign_d;
  assign ifm_dff_x_12_11 = uSystolicPE_429_io_ifm_dff_d;
  assign uSystolicPE_429_io_enable_w = enable_w_x_10[12];
  assign uSystolicPE_429_io_clear_w = clear_w_x_10[12];
  assign wght_sign_x_10_13 = uSystolicPE_429_io_wght_sign_d;
  assign wght_abs_x_10_13 = uSystolicPE_429_io_wght_abs_d;
  assign uSystolicPE_429_io_enable_o = enable_o_x_10[13];
  assign uSystolicPE_429_io_clear_o = clear_o_x_10[13];
  assign ofm_x_10_12 = uSystolicPE_429_io_ofm_d;
  assign randW_x_12_11 = uSystolicPE_429_io_randW_d;
  assign uSystolicPE_430_io_mac_done = mac_done_x_12[11];
  assign uSystolicPE_430_io_enable_i = enable_i_x_12[11];
  assign uSystolicPE_430_io_clear_i = clear_i_x_12[11];
  assign ifm_sign_x_12_12 = uSystolicPE_430_io_ifm_sign_d;
  assign ifm_dff_x_12_12 = uSystolicPE_430_io_ifm_dff_d;
  assign uSystolicPE_430_io_enable_w = enable_w_x_11[12];
  assign uSystolicPE_430_io_clear_w = clear_w_x_11[12];
  assign wght_sign_x_11_13 = uSystolicPE_430_io_wght_sign_d;
  assign wght_abs_x_11_13 = uSystolicPE_430_io_wght_abs_d;
  assign uSystolicPE_430_io_enable_o = enable_o_x_11[13];
  assign uSystolicPE_430_io_clear_o = clear_o_x_11[13];
  assign ofm_x_11_12 = uSystolicPE_430_io_ofm_d;
  assign randW_x_12_12 = uSystolicPE_430_io_randW_d;
  assign uSystolicPE_431_io_mac_done = mac_done_x_12[12];
  assign uSystolicPE_431_io_enable_i = enable_i_x_12[12];
  assign uSystolicPE_431_io_clear_i = clear_i_x_12[12];
  assign ifm_sign_x_12_13 = uSystolicPE_431_io_ifm_sign_d;
  assign ifm_dff_x_12_13 = uSystolicPE_431_io_ifm_dff_d;
  assign uSystolicPE_431_io_enable_w = enable_w_x_12[12];
  assign uSystolicPE_431_io_clear_w = clear_w_x_12[12];
  assign wght_sign_x_12_13 = uSystolicPE_431_io_wght_sign_d;
  assign wght_abs_x_12_13 = uSystolicPE_431_io_wght_abs_d;
  assign uSystolicPE_431_io_enable_o = enable_o_x_12[13];
  assign uSystolicPE_431_io_clear_o = clear_o_x_12[13];
  assign ofm_x_12_12 = uSystolicPE_431_io_ofm_d;
  assign randW_x_12_13 = uSystolicPE_431_io_randW_d;
  assign uSystolicPE_432_io_mac_done = mac_done_x_12[13];
  assign uSystolicPE_432_io_enable_i = enable_i_x_12[13];
  assign uSystolicPE_432_io_clear_i = clear_i_x_12[13];
  assign ifm_sign_x_12_14 = uSystolicPE_432_io_ifm_sign_d;
  assign ifm_dff_x_12_14 = uSystolicPE_432_io_ifm_dff_d;
  assign uSystolicPE_432_io_enable_w = enable_w_x_13[12];
  assign uSystolicPE_432_io_clear_w = clear_w_x_13[12];
  assign wght_sign_x_13_13 = uSystolicPE_432_io_wght_sign_d;
  assign wght_abs_x_13_13 = uSystolicPE_432_io_wght_abs_d;
  assign uSystolicPE_432_io_enable_o = enable_o_x_13[13];
  assign uSystolicPE_432_io_clear_o = clear_o_x_13[13];
  assign ofm_x_13_12 = uSystolicPE_432_io_ofm_d;
  assign randW_x_12_14 = uSystolicPE_432_io_randW_d;
  assign uSystolicPE_433_io_mac_done = mac_done_x_12[14];
  assign uSystolicPE_433_io_enable_i = enable_i_x_12[14];
  assign uSystolicPE_433_io_clear_i = clear_i_x_12[14];
  assign ifm_sign_x_12_15 = uSystolicPE_433_io_ifm_sign_d;
  assign ifm_dff_x_12_15 = uSystolicPE_433_io_ifm_dff_d;
  assign uSystolicPE_433_io_enable_w = enable_w_x_14[12];
  assign uSystolicPE_433_io_clear_w = clear_w_x_14[12];
  assign wght_sign_x_14_13 = uSystolicPE_433_io_wght_sign_d;
  assign wght_abs_x_14_13 = uSystolicPE_433_io_wght_abs_d;
  assign uSystolicPE_433_io_enable_o = enable_o_x_14[13];
  assign uSystolicPE_433_io_clear_o = clear_o_x_14[13];
  assign ofm_x_14_12 = uSystolicPE_433_io_ofm_d;
  assign randW_x_12_15 = uSystolicPE_433_io_randW_d;
  assign uSystolicPE_434_io_mac_done = mac_done_x_12[15];
  assign uSystolicPE_434_io_enable_i = enable_i_x_12[15];
  assign uSystolicPE_434_io_clear_i = clear_i_x_12[15];
  assign ifm_sign_x_12_16 = uSystolicPE_434_io_ifm_sign_d;
  assign ifm_dff_x_12_16 = uSystolicPE_434_io_ifm_dff_d;
  assign uSystolicPE_434_io_enable_w = enable_w_x_15[12];
  assign uSystolicPE_434_io_clear_w = clear_w_x_15[12];
  assign wght_sign_x_15_13 = uSystolicPE_434_io_wght_sign_d;
  assign wght_abs_x_15_13 = uSystolicPE_434_io_wght_abs_d;
  assign uSystolicPE_434_io_enable_o = enable_o_x_15[13];
  assign uSystolicPE_434_io_clear_o = clear_o_x_15[13];
  assign ofm_x_15_12 = uSystolicPE_434_io_ofm_d;
  assign randW_x_12_16 = uSystolicPE_434_io_randW_d;
  assign uSystolicPEBorder_29_io_mac_done = mac_done_x_13[0];
  assign uSystolicPEBorder_29_io_enable_i = enable_i_x_13[0];
  assign uSystolicPEBorder_29_io_clear_i = clear_i_x_13[0];
  assign ifm_sign_x_13_1 = uSystolicPEBorder_29_io_ifm_sign_d;
  assign ifm_dff_x_13_1 = uSystolicPEBorder_29_io_ifm_dff_d;
  assign uSystolicPEBorder_29_io_enable_w = enable_w_x_0[13];
  assign uSystolicPEBorder_29_io_clear_w = clear_w_x_0[13];
  assign wght_sign_x_0_14 = uSystolicPEBorder_29_io_wght_sign_d;
  assign wght_abs_x_0_14 = uSystolicPEBorder_29_io_wght_abs_d;
  assign uSystolicPEBorder_29_io_enable_o = enable_o_x_0[14];
  assign uSystolicPEBorder_29_io_clear_o = clear_o_x_0[14];
  assign ofm_x_0_13 = uSystolicPEBorder_29_io_ofm_d;
  assign randW_x_13_1 = uSystolicPEBorder_29_io_randW_d;
  assign uSystolicPE_435_io_mac_done = mac_done_x_13[1];
  assign uSystolicPE_435_io_enable_i = enable_i_x_13[1];
  assign uSystolicPE_435_io_clear_i = clear_i_x_13[1];
  assign ifm_sign_x_13_2 = uSystolicPE_435_io_ifm_sign_d;
  assign ifm_dff_x_13_2 = uSystolicPE_435_io_ifm_dff_d;
  assign uSystolicPE_435_io_enable_w = enable_w_x_1[13];
  assign uSystolicPE_435_io_clear_w = clear_w_x_1[13];
  assign wght_sign_x_1_14 = uSystolicPE_435_io_wght_sign_d;
  assign wght_abs_x_1_14 = uSystolicPE_435_io_wght_abs_d;
  assign uSystolicPE_435_io_enable_o = enable_o_x_1[14];
  assign uSystolicPE_435_io_clear_o = clear_o_x_1[14];
  assign ofm_x_1_13 = uSystolicPE_435_io_ofm_d;
  assign randW_x_13_2 = uSystolicPE_435_io_randW_d;
  assign uSystolicPE_436_io_mac_done = mac_done_x_13[2];
  assign uSystolicPE_436_io_enable_i = enable_i_x_13[2];
  assign uSystolicPE_436_io_clear_i = clear_i_x_13[2];
  assign ifm_sign_x_13_3 = uSystolicPE_436_io_ifm_sign_d;
  assign ifm_dff_x_13_3 = uSystolicPE_436_io_ifm_dff_d;
  assign uSystolicPE_436_io_enable_w = enable_w_x_2[13];
  assign uSystolicPE_436_io_clear_w = clear_w_x_2[13];
  assign wght_sign_x_2_14 = uSystolicPE_436_io_wght_sign_d;
  assign wght_abs_x_2_14 = uSystolicPE_436_io_wght_abs_d;
  assign uSystolicPE_436_io_enable_o = enable_o_x_2[14];
  assign uSystolicPE_436_io_clear_o = clear_o_x_2[14];
  assign ofm_x_2_13 = uSystolicPE_436_io_ofm_d;
  assign randW_x_13_3 = uSystolicPE_436_io_randW_d;
  assign uSystolicPE_437_io_mac_done = mac_done_x_13[3];
  assign uSystolicPE_437_io_enable_i = enable_i_x_13[3];
  assign uSystolicPE_437_io_clear_i = clear_i_x_13[3];
  assign ifm_sign_x_13_4 = uSystolicPE_437_io_ifm_sign_d;
  assign ifm_dff_x_13_4 = uSystolicPE_437_io_ifm_dff_d;
  assign uSystolicPE_437_io_enable_w = enable_w_x_3[13];
  assign uSystolicPE_437_io_clear_w = clear_w_x_3[13];
  assign wght_sign_x_3_14 = uSystolicPE_437_io_wght_sign_d;
  assign wght_abs_x_3_14 = uSystolicPE_437_io_wght_abs_d;
  assign uSystolicPE_437_io_enable_o = enable_o_x_3[14];
  assign uSystolicPE_437_io_clear_o = clear_o_x_3[14];
  assign ofm_x_3_13 = uSystolicPE_437_io_ofm_d;
  assign randW_x_13_4 = uSystolicPE_437_io_randW_d;
  assign uSystolicPE_438_io_mac_done = mac_done_x_13[4];
  assign uSystolicPE_438_io_enable_i = enable_i_x_13[4];
  assign uSystolicPE_438_io_clear_i = clear_i_x_13[4];
  assign ifm_sign_x_13_5 = uSystolicPE_438_io_ifm_sign_d;
  assign ifm_dff_x_13_5 = uSystolicPE_438_io_ifm_dff_d;
  assign uSystolicPE_438_io_enable_w = enable_w_x_4[13];
  assign uSystolicPE_438_io_clear_w = clear_w_x_4[13];
  assign wght_sign_x_4_14 = uSystolicPE_438_io_wght_sign_d;
  assign wght_abs_x_4_14 = uSystolicPE_438_io_wght_abs_d;
  assign uSystolicPE_438_io_enable_o = enable_o_x_4[14];
  assign uSystolicPE_438_io_clear_o = clear_o_x_4[14];
  assign ofm_x_4_13 = uSystolicPE_438_io_ofm_d;
  assign randW_x_13_5 = uSystolicPE_438_io_randW_d;
  assign uSystolicPE_439_io_mac_done = mac_done_x_13[5];
  assign uSystolicPE_439_io_enable_i = enable_i_x_13[5];
  assign uSystolicPE_439_io_clear_i = clear_i_x_13[5];
  assign ifm_sign_x_13_6 = uSystolicPE_439_io_ifm_sign_d;
  assign ifm_dff_x_13_6 = uSystolicPE_439_io_ifm_dff_d;
  assign uSystolicPE_439_io_enable_w = enable_w_x_5[13];
  assign uSystolicPE_439_io_clear_w = clear_w_x_5[13];
  assign wght_sign_x_5_14 = uSystolicPE_439_io_wght_sign_d;
  assign wght_abs_x_5_14 = uSystolicPE_439_io_wght_abs_d;
  assign uSystolicPE_439_io_enable_o = enable_o_x_5[14];
  assign uSystolicPE_439_io_clear_o = clear_o_x_5[14];
  assign ofm_x_5_13 = uSystolicPE_439_io_ofm_d;
  assign randW_x_13_6 = uSystolicPE_439_io_randW_d;
  assign uSystolicPE_440_io_mac_done = mac_done_x_13[6];
  assign uSystolicPE_440_io_enable_i = enable_i_x_13[6];
  assign uSystolicPE_440_io_clear_i = clear_i_x_13[6];
  assign ifm_sign_x_13_7 = uSystolicPE_440_io_ifm_sign_d;
  assign ifm_dff_x_13_7 = uSystolicPE_440_io_ifm_dff_d;
  assign uSystolicPE_440_io_enable_w = enable_w_x_6[13];
  assign uSystolicPE_440_io_clear_w = clear_w_x_6[13];
  assign wght_sign_x_6_14 = uSystolicPE_440_io_wght_sign_d;
  assign wght_abs_x_6_14 = uSystolicPE_440_io_wght_abs_d;
  assign uSystolicPE_440_io_enable_o = enable_o_x_6[14];
  assign uSystolicPE_440_io_clear_o = clear_o_x_6[14];
  assign ofm_x_6_13 = uSystolicPE_440_io_ofm_d;
  assign randW_x_13_7 = uSystolicPE_440_io_randW_d;
  assign uSystolicPE_441_io_mac_done = mac_done_x_13[7];
  assign uSystolicPE_441_io_enable_i = enable_i_x_13[7];
  assign uSystolicPE_441_io_clear_i = clear_i_x_13[7];
  assign ifm_sign_x_13_8 = uSystolicPE_441_io_ifm_sign_d;
  assign ifm_dff_x_13_8 = uSystolicPE_441_io_ifm_dff_d;
  assign uSystolicPE_441_io_enable_w = enable_w_x_7[13];
  assign uSystolicPE_441_io_clear_w = clear_w_x_7[13];
  assign wght_sign_x_7_14 = uSystolicPE_441_io_wght_sign_d;
  assign wght_abs_x_7_14 = uSystolicPE_441_io_wght_abs_d;
  assign uSystolicPE_441_io_enable_o = enable_o_x_7[14];
  assign uSystolicPE_441_io_clear_o = clear_o_x_7[14];
  assign ofm_x_7_13 = uSystolicPE_441_io_ofm_d;
  assign randW_x_13_8 = uSystolicPE_441_io_randW_d;
  assign uSystolicPE_442_io_mac_done = mac_done_x_13[8];
  assign uSystolicPE_442_io_enable_i = enable_i_x_13[8];
  assign uSystolicPE_442_io_clear_i = clear_i_x_13[8];
  assign ifm_sign_x_13_9 = uSystolicPE_442_io_ifm_sign_d;
  assign ifm_dff_x_13_9 = uSystolicPE_442_io_ifm_dff_d;
  assign uSystolicPE_442_io_enable_w = enable_w_x_8[13];
  assign uSystolicPE_442_io_clear_w = clear_w_x_8[13];
  assign wght_sign_x_8_14 = uSystolicPE_442_io_wght_sign_d;
  assign wght_abs_x_8_14 = uSystolicPE_442_io_wght_abs_d;
  assign uSystolicPE_442_io_enable_o = enable_o_x_8[14];
  assign uSystolicPE_442_io_clear_o = clear_o_x_8[14];
  assign ofm_x_8_13 = uSystolicPE_442_io_ofm_d;
  assign randW_x_13_9 = uSystolicPE_442_io_randW_d;
  assign uSystolicPE_443_io_mac_done = mac_done_x_13[9];
  assign uSystolicPE_443_io_enable_i = enable_i_x_13[9];
  assign uSystolicPE_443_io_clear_i = clear_i_x_13[9];
  assign ifm_sign_x_13_10 = uSystolicPE_443_io_ifm_sign_d;
  assign ifm_dff_x_13_10 = uSystolicPE_443_io_ifm_dff_d;
  assign uSystolicPE_443_io_enable_w = enable_w_x_9[13];
  assign uSystolicPE_443_io_clear_w = clear_w_x_9[13];
  assign wght_sign_x_9_14 = uSystolicPE_443_io_wght_sign_d;
  assign wght_abs_x_9_14 = uSystolicPE_443_io_wght_abs_d;
  assign uSystolicPE_443_io_enable_o = enable_o_x_9[14];
  assign uSystolicPE_443_io_clear_o = clear_o_x_9[14];
  assign ofm_x_9_13 = uSystolicPE_443_io_ofm_d;
  assign randW_x_13_10 = uSystolicPE_443_io_randW_d;
  assign uSystolicPE_444_io_mac_done = mac_done_x_13[10];
  assign uSystolicPE_444_io_enable_i = enable_i_x_13[10];
  assign uSystolicPE_444_io_clear_i = clear_i_x_13[10];
  assign ifm_sign_x_13_11 = uSystolicPE_444_io_ifm_sign_d;
  assign ifm_dff_x_13_11 = uSystolicPE_444_io_ifm_dff_d;
  assign uSystolicPE_444_io_enable_w = enable_w_x_10[13];
  assign uSystolicPE_444_io_clear_w = clear_w_x_10[13];
  assign wght_sign_x_10_14 = uSystolicPE_444_io_wght_sign_d;
  assign wght_abs_x_10_14 = uSystolicPE_444_io_wght_abs_d;
  assign uSystolicPE_444_io_enable_o = enable_o_x_10[14];
  assign uSystolicPE_444_io_clear_o = clear_o_x_10[14];
  assign ofm_x_10_13 = uSystolicPE_444_io_ofm_d;
  assign randW_x_13_11 = uSystolicPE_444_io_randW_d;
  assign uSystolicPE_445_io_mac_done = mac_done_x_13[11];
  assign uSystolicPE_445_io_enable_i = enable_i_x_13[11];
  assign uSystolicPE_445_io_clear_i = clear_i_x_13[11];
  assign ifm_sign_x_13_12 = uSystolicPE_445_io_ifm_sign_d;
  assign ifm_dff_x_13_12 = uSystolicPE_445_io_ifm_dff_d;
  assign uSystolicPE_445_io_enable_w = enable_w_x_11[13];
  assign uSystolicPE_445_io_clear_w = clear_w_x_11[13];
  assign wght_sign_x_11_14 = uSystolicPE_445_io_wght_sign_d;
  assign wght_abs_x_11_14 = uSystolicPE_445_io_wght_abs_d;
  assign uSystolicPE_445_io_enable_o = enable_o_x_11[14];
  assign uSystolicPE_445_io_clear_o = clear_o_x_11[14];
  assign ofm_x_11_13 = uSystolicPE_445_io_ofm_d;
  assign randW_x_13_12 = uSystolicPE_445_io_randW_d;
  assign uSystolicPE_446_io_mac_done = mac_done_x_13[12];
  assign uSystolicPE_446_io_enable_i = enable_i_x_13[12];
  assign uSystolicPE_446_io_clear_i = clear_i_x_13[12];
  assign ifm_sign_x_13_13 = uSystolicPE_446_io_ifm_sign_d;
  assign ifm_dff_x_13_13 = uSystolicPE_446_io_ifm_dff_d;
  assign uSystolicPE_446_io_enable_w = enable_w_x_12[13];
  assign uSystolicPE_446_io_clear_w = clear_w_x_12[13];
  assign wght_sign_x_12_14 = uSystolicPE_446_io_wght_sign_d;
  assign wght_abs_x_12_14 = uSystolicPE_446_io_wght_abs_d;
  assign uSystolicPE_446_io_enable_o = enable_o_x_12[14];
  assign uSystolicPE_446_io_clear_o = clear_o_x_12[14];
  assign ofm_x_12_13 = uSystolicPE_446_io_ofm_d;
  assign randW_x_13_13 = uSystolicPE_446_io_randW_d;
  assign uSystolicPE_447_io_mac_done = mac_done_x_13[13];
  assign uSystolicPE_447_io_enable_i = enable_i_x_13[13];
  assign uSystolicPE_447_io_clear_i = clear_i_x_13[13];
  assign ifm_sign_x_13_14 = uSystolicPE_447_io_ifm_sign_d;
  assign ifm_dff_x_13_14 = uSystolicPE_447_io_ifm_dff_d;
  assign uSystolicPE_447_io_enable_w = enable_w_x_13[13];
  assign uSystolicPE_447_io_clear_w = clear_w_x_13[13];
  assign wght_sign_x_13_14 = uSystolicPE_447_io_wght_sign_d;
  assign wght_abs_x_13_14 = uSystolicPE_447_io_wght_abs_d;
  assign uSystolicPE_447_io_enable_o = enable_o_x_13[14];
  assign uSystolicPE_447_io_clear_o = clear_o_x_13[14];
  assign ofm_x_13_13 = uSystolicPE_447_io_ofm_d;
  assign randW_x_13_14 = uSystolicPE_447_io_randW_d;
  assign uSystolicPE_448_io_mac_done = mac_done_x_13[14];
  assign uSystolicPE_448_io_enable_i = enable_i_x_13[14];
  assign uSystolicPE_448_io_clear_i = clear_i_x_13[14];
  assign ifm_sign_x_13_15 = uSystolicPE_448_io_ifm_sign_d;
  assign ifm_dff_x_13_15 = uSystolicPE_448_io_ifm_dff_d;
  assign uSystolicPE_448_io_enable_w = enable_w_x_14[13];
  assign uSystolicPE_448_io_clear_w = clear_w_x_14[13];
  assign wght_sign_x_14_14 = uSystolicPE_448_io_wght_sign_d;
  assign wght_abs_x_14_14 = uSystolicPE_448_io_wght_abs_d;
  assign uSystolicPE_448_io_enable_o = enable_o_x_14[14];
  assign uSystolicPE_448_io_clear_o = clear_o_x_14[14];
  assign ofm_x_14_13 = uSystolicPE_448_io_ofm_d;
  assign randW_x_13_15 = uSystolicPE_448_io_randW_d;
  assign uSystolicPE_449_io_mac_done = mac_done_x_13[15];
  assign uSystolicPE_449_io_enable_i = enable_i_x_13[15];
  assign uSystolicPE_449_io_clear_i = clear_i_x_13[15];
  assign ifm_sign_x_13_16 = uSystolicPE_449_io_ifm_sign_d;
  assign ifm_dff_x_13_16 = uSystolicPE_449_io_ifm_dff_d;
  assign uSystolicPE_449_io_enable_w = enable_w_x_15[13];
  assign uSystolicPE_449_io_clear_w = clear_w_x_15[13];
  assign wght_sign_x_15_14 = uSystolicPE_449_io_wght_sign_d;
  assign wght_abs_x_15_14 = uSystolicPE_449_io_wght_abs_d;
  assign uSystolicPE_449_io_enable_o = enable_o_x_15[14];
  assign uSystolicPE_449_io_clear_o = clear_o_x_15[14];
  assign ofm_x_15_13 = uSystolicPE_449_io_ofm_d;
  assign randW_x_13_16 = uSystolicPE_449_io_randW_d;
  assign uSystolicPEBorder_30_io_mac_done = mac_done_x_14[0];
  assign uSystolicPEBorder_30_io_enable_i = enable_i_x_14[0];
  assign uSystolicPEBorder_30_io_clear_i = clear_i_x_14[0];
  assign ifm_sign_x_14_1 = uSystolicPEBorder_30_io_ifm_sign_d;
  assign ifm_dff_x_14_1 = uSystolicPEBorder_30_io_ifm_dff_d;
  assign uSystolicPEBorder_30_io_enable_w = enable_w_x_0[14];
  assign uSystolicPEBorder_30_io_clear_w = clear_w_x_0[14];
  assign wght_sign_x_0_15 = uSystolicPEBorder_30_io_wght_sign_d;
  assign wght_abs_x_0_15 = uSystolicPEBorder_30_io_wght_abs_d;
  assign uSystolicPEBorder_30_io_enable_o = enable_o_x_0[15];
  assign uSystolicPEBorder_30_io_clear_o = clear_o_x_0[15];
  assign ofm_x_0_14 = uSystolicPEBorder_30_io_ofm_d;
  assign randW_x_14_1 = uSystolicPEBorder_30_io_randW_d;
  assign uSystolicPE_450_io_mac_done = mac_done_x_14[1];
  assign uSystolicPE_450_io_enable_i = enable_i_x_14[1];
  assign uSystolicPE_450_io_clear_i = clear_i_x_14[1];
  assign ifm_sign_x_14_2 = uSystolicPE_450_io_ifm_sign_d;
  assign ifm_dff_x_14_2 = uSystolicPE_450_io_ifm_dff_d;
  assign uSystolicPE_450_io_enable_w = enable_w_x_1[14];
  assign uSystolicPE_450_io_clear_w = clear_w_x_1[14];
  assign wght_sign_x_1_15 = uSystolicPE_450_io_wght_sign_d;
  assign wght_abs_x_1_15 = uSystolicPE_450_io_wght_abs_d;
  assign uSystolicPE_450_io_enable_o = enable_o_x_1[15];
  assign uSystolicPE_450_io_clear_o = clear_o_x_1[15];
  assign ofm_x_1_14 = uSystolicPE_450_io_ofm_d;
  assign randW_x_14_2 = uSystolicPE_450_io_randW_d;
  assign uSystolicPE_451_io_mac_done = mac_done_x_14[2];
  assign uSystolicPE_451_io_enable_i = enable_i_x_14[2];
  assign uSystolicPE_451_io_clear_i = clear_i_x_14[2];
  assign ifm_sign_x_14_3 = uSystolicPE_451_io_ifm_sign_d;
  assign ifm_dff_x_14_3 = uSystolicPE_451_io_ifm_dff_d;
  assign uSystolicPE_451_io_enable_w = enable_w_x_2[14];
  assign uSystolicPE_451_io_clear_w = clear_w_x_2[14];
  assign wght_sign_x_2_15 = uSystolicPE_451_io_wght_sign_d;
  assign wght_abs_x_2_15 = uSystolicPE_451_io_wght_abs_d;
  assign uSystolicPE_451_io_enable_o = enable_o_x_2[15];
  assign uSystolicPE_451_io_clear_o = clear_o_x_2[15];
  assign ofm_x_2_14 = uSystolicPE_451_io_ofm_d;
  assign randW_x_14_3 = uSystolicPE_451_io_randW_d;
  assign uSystolicPE_452_io_mac_done = mac_done_x_14[3];
  assign uSystolicPE_452_io_enable_i = enable_i_x_14[3];
  assign uSystolicPE_452_io_clear_i = clear_i_x_14[3];
  assign ifm_sign_x_14_4 = uSystolicPE_452_io_ifm_sign_d;
  assign ifm_dff_x_14_4 = uSystolicPE_452_io_ifm_dff_d;
  assign uSystolicPE_452_io_enable_w = enable_w_x_3[14];
  assign uSystolicPE_452_io_clear_w = clear_w_x_3[14];
  assign wght_sign_x_3_15 = uSystolicPE_452_io_wght_sign_d;
  assign wght_abs_x_3_15 = uSystolicPE_452_io_wght_abs_d;
  assign uSystolicPE_452_io_enable_o = enable_o_x_3[15];
  assign uSystolicPE_452_io_clear_o = clear_o_x_3[15];
  assign ofm_x_3_14 = uSystolicPE_452_io_ofm_d;
  assign randW_x_14_4 = uSystolicPE_452_io_randW_d;
  assign uSystolicPE_453_io_mac_done = mac_done_x_14[4];
  assign uSystolicPE_453_io_enable_i = enable_i_x_14[4];
  assign uSystolicPE_453_io_clear_i = clear_i_x_14[4];
  assign ifm_sign_x_14_5 = uSystolicPE_453_io_ifm_sign_d;
  assign ifm_dff_x_14_5 = uSystolicPE_453_io_ifm_dff_d;
  assign uSystolicPE_453_io_enable_w = enable_w_x_4[14];
  assign uSystolicPE_453_io_clear_w = clear_w_x_4[14];
  assign wght_sign_x_4_15 = uSystolicPE_453_io_wght_sign_d;
  assign wght_abs_x_4_15 = uSystolicPE_453_io_wght_abs_d;
  assign uSystolicPE_453_io_enable_o = enable_o_x_4[15];
  assign uSystolicPE_453_io_clear_o = clear_o_x_4[15];
  assign ofm_x_4_14 = uSystolicPE_453_io_ofm_d;
  assign randW_x_14_5 = uSystolicPE_453_io_randW_d;
  assign uSystolicPE_454_io_mac_done = mac_done_x_14[5];
  assign uSystolicPE_454_io_enable_i = enable_i_x_14[5];
  assign uSystolicPE_454_io_clear_i = clear_i_x_14[5];
  assign ifm_sign_x_14_6 = uSystolicPE_454_io_ifm_sign_d;
  assign ifm_dff_x_14_6 = uSystolicPE_454_io_ifm_dff_d;
  assign uSystolicPE_454_io_enable_w = enable_w_x_5[14];
  assign uSystolicPE_454_io_clear_w = clear_w_x_5[14];
  assign wght_sign_x_5_15 = uSystolicPE_454_io_wght_sign_d;
  assign wght_abs_x_5_15 = uSystolicPE_454_io_wght_abs_d;
  assign uSystolicPE_454_io_enable_o = enable_o_x_5[15];
  assign uSystolicPE_454_io_clear_o = clear_o_x_5[15];
  assign ofm_x_5_14 = uSystolicPE_454_io_ofm_d;
  assign randW_x_14_6 = uSystolicPE_454_io_randW_d;
  assign uSystolicPE_455_io_mac_done = mac_done_x_14[6];
  assign uSystolicPE_455_io_enable_i = enable_i_x_14[6];
  assign uSystolicPE_455_io_clear_i = clear_i_x_14[6];
  assign ifm_sign_x_14_7 = uSystolicPE_455_io_ifm_sign_d;
  assign ifm_dff_x_14_7 = uSystolicPE_455_io_ifm_dff_d;
  assign uSystolicPE_455_io_enable_w = enable_w_x_6[14];
  assign uSystolicPE_455_io_clear_w = clear_w_x_6[14];
  assign wght_sign_x_6_15 = uSystolicPE_455_io_wght_sign_d;
  assign wght_abs_x_6_15 = uSystolicPE_455_io_wght_abs_d;
  assign uSystolicPE_455_io_enable_o = enable_o_x_6[15];
  assign uSystolicPE_455_io_clear_o = clear_o_x_6[15];
  assign ofm_x_6_14 = uSystolicPE_455_io_ofm_d;
  assign randW_x_14_7 = uSystolicPE_455_io_randW_d;
  assign uSystolicPE_456_io_mac_done = mac_done_x_14[7];
  assign uSystolicPE_456_io_enable_i = enable_i_x_14[7];
  assign uSystolicPE_456_io_clear_i = clear_i_x_14[7];
  assign ifm_sign_x_14_8 = uSystolicPE_456_io_ifm_sign_d;
  assign ifm_dff_x_14_8 = uSystolicPE_456_io_ifm_dff_d;
  assign uSystolicPE_456_io_enable_w = enable_w_x_7[14];
  assign uSystolicPE_456_io_clear_w = clear_w_x_7[14];
  assign wght_sign_x_7_15 = uSystolicPE_456_io_wght_sign_d;
  assign wght_abs_x_7_15 = uSystolicPE_456_io_wght_abs_d;
  assign uSystolicPE_456_io_enable_o = enable_o_x_7[15];
  assign uSystolicPE_456_io_clear_o = clear_o_x_7[15];
  assign ofm_x_7_14 = uSystolicPE_456_io_ofm_d;
  assign randW_x_14_8 = uSystolicPE_456_io_randW_d;
  assign uSystolicPE_457_io_mac_done = mac_done_x_14[8];
  assign uSystolicPE_457_io_enable_i = enable_i_x_14[8];
  assign uSystolicPE_457_io_clear_i = clear_i_x_14[8];
  assign ifm_sign_x_14_9 = uSystolicPE_457_io_ifm_sign_d;
  assign ifm_dff_x_14_9 = uSystolicPE_457_io_ifm_dff_d;
  assign uSystolicPE_457_io_enable_w = enable_w_x_8[14];
  assign uSystolicPE_457_io_clear_w = clear_w_x_8[14];
  assign wght_sign_x_8_15 = uSystolicPE_457_io_wght_sign_d;
  assign wght_abs_x_8_15 = uSystolicPE_457_io_wght_abs_d;
  assign uSystolicPE_457_io_enable_o = enable_o_x_8[15];
  assign uSystolicPE_457_io_clear_o = clear_o_x_8[15];
  assign ofm_x_8_14 = uSystolicPE_457_io_ofm_d;
  assign randW_x_14_9 = uSystolicPE_457_io_randW_d;
  assign uSystolicPE_458_io_mac_done = mac_done_x_14[9];
  assign uSystolicPE_458_io_enable_i = enable_i_x_14[9];
  assign uSystolicPE_458_io_clear_i = clear_i_x_14[9];
  assign ifm_sign_x_14_10 = uSystolicPE_458_io_ifm_sign_d;
  assign ifm_dff_x_14_10 = uSystolicPE_458_io_ifm_dff_d;
  assign uSystolicPE_458_io_enable_w = enable_w_x_9[14];
  assign uSystolicPE_458_io_clear_w = clear_w_x_9[14];
  assign wght_sign_x_9_15 = uSystolicPE_458_io_wght_sign_d;
  assign wght_abs_x_9_15 = uSystolicPE_458_io_wght_abs_d;
  assign uSystolicPE_458_io_enable_o = enable_o_x_9[15];
  assign uSystolicPE_458_io_clear_o = clear_o_x_9[15];
  assign ofm_x_9_14 = uSystolicPE_458_io_ofm_d;
  assign randW_x_14_10 = uSystolicPE_458_io_randW_d;
  assign uSystolicPE_459_io_mac_done = mac_done_x_14[10];
  assign uSystolicPE_459_io_enable_i = enable_i_x_14[10];
  assign uSystolicPE_459_io_clear_i = clear_i_x_14[10];
  assign ifm_sign_x_14_11 = uSystolicPE_459_io_ifm_sign_d;
  assign ifm_dff_x_14_11 = uSystolicPE_459_io_ifm_dff_d;
  assign uSystolicPE_459_io_enable_w = enable_w_x_10[14];
  assign uSystolicPE_459_io_clear_w = clear_w_x_10[14];
  assign wght_sign_x_10_15 = uSystolicPE_459_io_wght_sign_d;
  assign wght_abs_x_10_15 = uSystolicPE_459_io_wght_abs_d;
  assign uSystolicPE_459_io_enable_o = enable_o_x_10[15];
  assign uSystolicPE_459_io_clear_o = clear_o_x_10[15];
  assign ofm_x_10_14 = uSystolicPE_459_io_ofm_d;
  assign randW_x_14_11 = uSystolicPE_459_io_randW_d;
  assign uSystolicPE_460_io_mac_done = mac_done_x_14[11];
  assign uSystolicPE_460_io_enable_i = enable_i_x_14[11];
  assign uSystolicPE_460_io_clear_i = clear_i_x_14[11];
  assign ifm_sign_x_14_12 = uSystolicPE_460_io_ifm_sign_d;
  assign ifm_dff_x_14_12 = uSystolicPE_460_io_ifm_dff_d;
  assign uSystolicPE_460_io_enable_w = enable_w_x_11[14];
  assign uSystolicPE_460_io_clear_w = clear_w_x_11[14];
  assign wght_sign_x_11_15 = uSystolicPE_460_io_wght_sign_d;
  assign wght_abs_x_11_15 = uSystolicPE_460_io_wght_abs_d;
  assign uSystolicPE_460_io_enable_o = enable_o_x_11[15];
  assign uSystolicPE_460_io_clear_o = clear_o_x_11[15];
  assign ofm_x_11_14 = uSystolicPE_460_io_ofm_d;
  assign randW_x_14_12 = uSystolicPE_460_io_randW_d;
  assign uSystolicPE_461_io_mac_done = mac_done_x_14[12];
  assign uSystolicPE_461_io_enable_i = enable_i_x_14[12];
  assign uSystolicPE_461_io_clear_i = clear_i_x_14[12];
  assign ifm_sign_x_14_13 = uSystolicPE_461_io_ifm_sign_d;
  assign ifm_dff_x_14_13 = uSystolicPE_461_io_ifm_dff_d;
  assign uSystolicPE_461_io_enable_w = enable_w_x_12[14];
  assign uSystolicPE_461_io_clear_w = clear_w_x_12[14];
  assign wght_sign_x_12_15 = uSystolicPE_461_io_wght_sign_d;
  assign wght_abs_x_12_15 = uSystolicPE_461_io_wght_abs_d;
  assign uSystolicPE_461_io_enable_o = enable_o_x_12[15];
  assign uSystolicPE_461_io_clear_o = clear_o_x_12[15];
  assign ofm_x_12_14 = uSystolicPE_461_io_ofm_d;
  assign randW_x_14_13 = uSystolicPE_461_io_randW_d;
  assign uSystolicPE_462_io_mac_done = mac_done_x_14[13];
  assign uSystolicPE_462_io_enable_i = enable_i_x_14[13];
  assign uSystolicPE_462_io_clear_i = clear_i_x_14[13];
  assign ifm_sign_x_14_14 = uSystolicPE_462_io_ifm_sign_d;
  assign ifm_dff_x_14_14 = uSystolicPE_462_io_ifm_dff_d;
  assign uSystolicPE_462_io_enable_w = enable_w_x_13[14];
  assign uSystolicPE_462_io_clear_w = clear_w_x_13[14];
  assign wght_sign_x_13_15 = uSystolicPE_462_io_wght_sign_d;
  assign wght_abs_x_13_15 = uSystolicPE_462_io_wght_abs_d;
  assign uSystolicPE_462_io_enable_o = enable_o_x_13[15];
  assign uSystolicPE_462_io_clear_o = clear_o_x_13[15];
  assign ofm_x_13_14 = uSystolicPE_462_io_ofm_d;
  assign randW_x_14_14 = uSystolicPE_462_io_randW_d;
  assign uSystolicPE_463_io_mac_done = mac_done_x_14[14];
  assign uSystolicPE_463_io_enable_i = enable_i_x_14[14];
  assign uSystolicPE_463_io_clear_i = clear_i_x_14[14];
  assign ifm_sign_x_14_15 = uSystolicPE_463_io_ifm_sign_d;
  assign ifm_dff_x_14_15 = uSystolicPE_463_io_ifm_dff_d;
  assign uSystolicPE_463_io_enable_w = enable_w_x_14[14];
  assign uSystolicPE_463_io_clear_w = clear_w_x_14[14];
  assign wght_sign_x_14_15 = uSystolicPE_463_io_wght_sign_d;
  assign wght_abs_x_14_15 = uSystolicPE_463_io_wght_abs_d;
  assign uSystolicPE_463_io_enable_o = enable_o_x_14[15];
  assign uSystolicPE_463_io_clear_o = clear_o_x_14[15];
  assign ofm_x_14_14 = uSystolicPE_463_io_ofm_d;
  assign randW_x_14_15 = uSystolicPE_463_io_randW_d;
  assign uSystolicPE_464_io_mac_done = mac_done_x_14[15];
  assign uSystolicPE_464_io_enable_i = enable_i_x_14[15];
  assign uSystolicPE_464_io_clear_i = clear_i_x_14[15];
  assign ifm_sign_x_14_16 = uSystolicPE_464_io_ifm_sign_d;
  assign ifm_dff_x_14_16 = uSystolicPE_464_io_ifm_dff_d;
  assign uSystolicPE_464_io_enable_w = enable_w_x_15[14];
  assign uSystolicPE_464_io_clear_w = clear_w_x_15[14];
  assign wght_sign_x_15_15 = uSystolicPE_464_io_wght_sign_d;
  assign wght_abs_x_15_15 = uSystolicPE_464_io_wght_abs_d;
  assign uSystolicPE_464_io_enable_o = enable_o_x_15[15];
  assign uSystolicPE_464_io_clear_o = clear_o_x_15[15];
  assign ofm_x_15_14 = uSystolicPE_464_io_ofm_d;
  assign randW_x_14_16 = uSystolicPE_464_io_randW_d;
  assign uSystolicPEBorder_31_io_mac_done = mac_done_x_15[0];
  assign uSystolicPEBorder_31_io_enable_i = enable_i_x_15[0];
  assign uSystolicPEBorder_31_io_clear_i = clear_i_x_15[0];
  assign ifm_sign_x_15_1 = uSystolicPEBorder_31_io_ifm_sign_d;
  assign ifm_dff_x_15_1 = uSystolicPEBorder_31_io_ifm_dff_d;
  assign uSystolicPEBorder_31_io_enable_w = enable_w_x_0[15];
  assign uSystolicPEBorder_31_io_clear_w = clear_w_x_0[15];
  assign wght_sign_x_0_16 = uSystolicPEBorder_31_io_wght_sign_d;
  assign wght_abs_x_0_16 = uSystolicPEBorder_31_io_wght_abs_d;
  assign uSystolicPEBorder_31_io_enable_o = enable_o_x_0[16];
  assign uSystolicPEBorder_31_io_clear_o = clear_o_x_0[16];
  assign ofm_x_0_15 = uSystolicPEBorder_31_io_ofm_d;
  assign randW_x_15_1 = uSystolicPEBorder_31_io_randW_d;
  assign uSystolicPE_465_io_mac_done = mac_done_x_15[1];
  assign uSystolicPE_465_io_enable_i = enable_i_x_15[1];
  assign uSystolicPE_465_io_clear_i = clear_i_x_15[1];
  assign ifm_sign_x_15_2 = uSystolicPE_465_io_ifm_sign_d;
  assign ifm_dff_x_15_2 = uSystolicPE_465_io_ifm_dff_d;
  assign uSystolicPE_465_io_enable_w = enable_w_x_1[15];
  assign uSystolicPE_465_io_clear_w = clear_w_x_1[15];
  assign wght_sign_x_1_16 = uSystolicPE_465_io_wght_sign_d;
  assign wght_abs_x_1_16 = uSystolicPE_465_io_wght_abs_d;
  assign uSystolicPE_465_io_enable_o = enable_o_x_1[16];
  assign uSystolicPE_465_io_clear_o = clear_o_x_1[16];
  assign ofm_x_1_15 = uSystolicPE_465_io_ofm_d;
  assign randW_x_15_2 = uSystolicPE_465_io_randW_d;
  assign uSystolicPE_466_io_mac_done = mac_done_x_15[2];
  assign uSystolicPE_466_io_enable_i = enable_i_x_15[2];
  assign uSystolicPE_466_io_clear_i = clear_i_x_15[2];
  assign ifm_sign_x_15_3 = uSystolicPE_466_io_ifm_sign_d;
  assign ifm_dff_x_15_3 = uSystolicPE_466_io_ifm_dff_d;
  assign uSystolicPE_466_io_enable_w = enable_w_x_2[15];
  assign uSystolicPE_466_io_clear_w = clear_w_x_2[15];
  assign wght_sign_x_2_16 = uSystolicPE_466_io_wght_sign_d;
  assign wght_abs_x_2_16 = uSystolicPE_466_io_wght_abs_d;
  assign uSystolicPE_466_io_enable_o = enable_o_x_2[16];
  assign uSystolicPE_466_io_clear_o = clear_o_x_2[16];
  assign ofm_x_2_15 = uSystolicPE_466_io_ofm_d;
  assign randW_x_15_3 = uSystolicPE_466_io_randW_d;
  assign uSystolicPE_467_io_mac_done = mac_done_x_15[3];
  assign uSystolicPE_467_io_enable_i = enable_i_x_15[3];
  assign uSystolicPE_467_io_clear_i = clear_i_x_15[3];
  assign ifm_sign_x_15_4 = uSystolicPE_467_io_ifm_sign_d;
  assign ifm_dff_x_15_4 = uSystolicPE_467_io_ifm_dff_d;
  assign uSystolicPE_467_io_enable_w = enable_w_x_3[15];
  assign uSystolicPE_467_io_clear_w = clear_w_x_3[15];
  assign wght_sign_x_3_16 = uSystolicPE_467_io_wght_sign_d;
  assign wght_abs_x_3_16 = uSystolicPE_467_io_wght_abs_d;
  assign uSystolicPE_467_io_enable_o = enable_o_x_3[16];
  assign uSystolicPE_467_io_clear_o = clear_o_x_3[16];
  assign ofm_x_3_15 = uSystolicPE_467_io_ofm_d;
  assign randW_x_15_4 = uSystolicPE_467_io_randW_d;
  assign uSystolicPE_468_io_mac_done = mac_done_x_15[4];
  assign uSystolicPE_468_io_enable_i = enable_i_x_15[4];
  assign uSystolicPE_468_io_clear_i = clear_i_x_15[4];
  assign ifm_sign_x_15_5 = uSystolicPE_468_io_ifm_sign_d;
  assign ifm_dff_x_15_5 = uSystolicPE_468_io_ifm_dff_d;
  assign uSystolicPE_468_io_enable_w = enable_w_x_4[15];
  assign uSystolicPE_468_io_clear_w = clear_w_x_4[15];
  assign wght_sign_x_4_16 = uSystolicPE_468_io_wght_sign_d;
  assign wght_abs_x_4_16 = uSystolicPE_468_io_wght_abs_d;
  assign uSystolicPE_468_io_enable_o = enable_o_x_4[16];
  assign uSystolicPE_468_io_clear_o = clear_o_x_4[16];
  assign ofm_x_4_15 = uSystolicPE_468_io_ofm_d;
  assign randW_x_15_5 = uSystolicPE_468_io_randW_d;
  assign uSystolicPE_469_io_mac_done = mac_done_x_15[5];
  assign uSystolicPE_469_io_enable_i = enable_i_x_15[5];
  assign uSystolicPE_469_io_clear_i = clear_i_x_15[5];
  assign ifm_sign_x_15_6 = uSystolicPE_469_io_ifm_sign_d;
  assign ifm_dff_x_15_6 = uSystolicPE_469_io_ifm_dff_d;
  assign uSystolicPE_469_io_enable_w = enable_w_x_5[15];
  assign uSystolicPE_469_io_clear_w = clear_w_x_5[15];
  assign wght_sign_x_5_16 = uSystolicPE_469_io_wght_sign_d;
  assign wght_abs_x_5_16 = uSystolicPE_469_io_wght_abs_d;
  assign uSystolicPE_469_io_enable_o = enable_o_x_5[16];
  assign uSystolicPE_469_io_clear_o = clear_o_x_5[16];
  assign ofm_x_5_15 = uSystolicPE_469_io_ofm_d;
  assign randW_x_15_6 = uSystolicPE_469_io_randW_d;
  assign uSystolicPE_470_io_mac_done = mac_done_x_15[6];
  assign uSystolicPE_470_io_enable_i = enable_i_x_15[6];
  assign uSystolicPE_470_io_clear_i = clear_i_x_15[6];
  assign ifm_sign_x_15_7 = uSystolicPE_470_io_ifm_sign_d;
  assign ifm_dff_x_15_7 = uSystolicPE_470_io_ifm_dff_d;
  assign uSystolicPE_470_io_enable_w = enable_w_x_6[15];
  assign uSystolicPE_470_io_clear_w = clear_w_x_6[15];
  assign wght_sign_x_6_16 = uSystolicPE_470_io_wght_sign_d;
  assign wght_abs_x_6_16 = uSystolicPE_470_io_wght_abs_d;
  assign uSystolicPE_470_io_enable_o = enable_o_x_6[16];
  assign uSystolicPE_470_io_clear_o = clear_o_x_6[16];
  assign ofm_x_6_15 = uSystolicPE_470_io_ofm_d;
  assign randW_x_15_7 = uSystolicPE_470_io_randW_d;
  assign uSystolicPE_471_io_mac_done = mac_done_x_15[7];
  assign uSystolicPE_471_io_enable_i = enable_i_x_15[7];
  assign uSystolicPE_471_io_clear_i = clear_i_x_15[7];
  assign ifm_sign_x_15_8 = uSystolicPE_471_io_ifm_sign_d;
  assign ifm_dff_x_15_8 = uSystolicPE_471_io_ifm_dff_d;
  assign uSystolicPE_471_io_enable_w = enable_w_x_7[15];
  assign uSystolicPE_471_io_clear_w = clear_w_x_7[15];
  assign wght_sign_x_7_16 = uSystolicPE_471_io_wght_sign_d;
  assign wght_abs_x_7_16 = uSystolicPE_471_io_wght_abs_d;
  assign uSystolicPE_471_io_enable_o = enable_o_x_7[16];
  assign uSystolicPE_471_io_clear_o = clear_o_x_7[16];
  assign ofm_x_7_15 = uSystolicPE_471_io_ofm_d;
  assign randW_x_15_8 = uSystolicPE_471_io_randW_d;
  assign uSystolicPE_472_io_mac_done = mac_done_x_15[8];
  assign uSystolicPE_472_io_enable_i = enable_i_x_15[8];
  assign uSystolicPE_472_io_clear_i = clear_i_x_15[8];
  assign ifm_sign_x_15_9 = uSystolicPE_472_io_ifm_sign_d;
  assign ifm_dff_x_15_9 = uSystolicPE_472_io_ifm_dff_d;
  assign uSystolicPE_472_io_enable_w = enable_w_x_8[15];
  assign uSystolicPE_472_io_clear_w = clear_w_x_8[15];
  assign wght_sign_x_8_16 = uSystolicPE_472_io_wght_sign_d;
  assign wght_abs_x_8_16 = uSystolicPE_472_io_wght_abs_d;
  assign uSystolicPE_472_io_enable_o = enable_o_x_8[16];
  assign uSystolicPE_472_io_clear_o = clear_o_x_8[16];
  assign ofm_x_8_15 = uSystolicPE_472_io_ofm_d;
  assign randW_x_15_9 = uSystolicPE_472_io_randW_d;
  assign uSystolicPE_473_io_mac_done = mac_done_x_15[9];
  assign uSystolicPE_473_io_enable_i = enable_i_x_15[9];
  assign uSystolicPE_473_io_clear_i = clear_i_x_15[9];
  assign ifm_sign_x_15_10 = uSystolicPE_473_io_ifm_sign_d;
  assign ifm_dff_x_15_10 = uSystolicPE_473_io_ifm_dff_d;
  assign uSystolicPE_473_io_enable_w = enable_w_x_9[15];
  assign uSystolicPE_473_io_clear_w = clear_w_x_9[15];
  assign wght_sign_x_9_16 = uSystolicPE_473_io_wght_sign_d;
  assign wght_abs_x_9_16 = uSystolicPE_473_io_wght_abs_d;
  assign uSystolicPE_473_io_enable_o = enable_o_x_9[16];
  assign uSystolicPE_473_io_clear_o = clear_o_x_9[16];
  assign ofm_x_9_15 = uSystolicPE_473_io_ofm_d;
  assign randW_x_15_10 = uSystolicPE_473_io_randW_d;
  assign uSystolicPE_474_io_mac_done = mac_done_x_15[10];
  assign uSystolicPE_474_io_enable_i = enable_i_x_15[10];
  assign uSystolicPE_474_io_clear_i = clear_i_x_15[10];
  assign ifm_sign_x_15_11 = uSystolicPE_474_io_ifm_sign_d;
  assign ifm_dff_x_15_11 = uSystolicPE_474_io_ifm_dff_d;
  assign uSystolicPE_474_io_enable_w = enable_w_x_10[15];
  assign uSystolicPE_474_io_clear_w = clear_w_x_10[15];
  assign wght_sign_x_10_16 = uSystolicPE_474_io_wght_sign_d;
  assign wght_abs_x_10_16 = uSystolicPE_474_io_wght_abs_d;
  assign uSystolicPE_474_io_enable_o = enable_o_x_10[16];
  assign uSystolicPE_474_io_clear_o = clear_o_x_10[16];
  assign ofm_x_10_15 = uSystolicPE_474_io_ofm_d;
  assign randW_x_15_11 = uSystolicPE_474_io_randW_d;
  assign uSystolicPE_475_io_mac_done = mac_done_x_15[11];
  assign uSystolicPE_475_io_enable_i = enable_i_x_15[11];
  assign uSystolicPE_475_io_clear_i = clear_i_x_15[11];
  assign ifm_sign_x_15_12 = uSystolicPE_475_io_ifm_sign_d;
  assign ifm_dff_x_15_12 = uSystolicPE_475_io_ifm_dff_d;
  assign uSystolicPE_475_io_enable_w = enable_w_x_11[15];
  assign uSystolicPE_475_io_clear_w = clear_w_x_11[15];
  assign wght_sign_x_11_16 = uSystolicPE_475_io_wght_sign_d;
  assign wght_abs_x_11_16 = uSystolicPE_475_io_wght_abs_d;
  assign uSystolicPE_475_io_enable_o = enable_o_x_11[16];
  assign uSystolicPE_475_io_clear_o = clear_o_x_11[16];
  assign ofm_x_11_15 = uSystolicPE_475_io_ofm_d;
  assign randW_x_15_12 = uSystolicPE_475_io_randW_d;
  assign uSystolicPE_476_io_mac_done = mac_done_x_15[12];
  assign uSystolicPE_476_io_enable_i = enable_i_x_15[12];
  assign uSystolicPE_476_io_clear_i = clear_i_x_15[12];
  assign ifm_sign_x_15_13 = uSystolicPE_476_io_ifm_sign_d;
  assign ifm_dff_x_15_13 = uSystolicPE_476_io_ifm_dff_d;
  assign uSystolicPE_476_io_enable_w = enable_w_x_12[15];
  assign uSystolicPE_476_io_clear_w = clear_w_x_12[15];
  assign wght_sign_x_12_16 = uSystolicPE_476_io_wght_sign_d;
  assign wght_abs_x_12_16 = uSystolicPE_476_io_wght_abs_d;
  assign uSystolicPE_476_io_enable_o = enable_o_x_12[16];
  assign uSystolicPE_476_io_clear_o = clear_o_x_12[16];
  assign ofm_x_12_15 = uSystolicPE_476_io_ofm_d;
  assign randW_x_15_13 = uSystolicPE_476_io_randW_d;
  assign uSystolicPE_477_io_mac_done = mac_done_x_15[13];
  assign uSystolicPE_477_io_enable_i = enable_i_x_15[13];
  assign uSystolicPE_477_io_clear_i = clear_i_x_15[13];
  assign ifm_sign_x_15_14 = uSystolicPE_477_io_ifm_sign_d;
  assign ifm_dff_x_15_14 = uSystolicPE_477_io_ifm_dff_d;
  assign uSystolicPE_477_io_enable_w = enable_w_x_13[15];
  assign uSystolicPE_477_io_clear_w = clear_w_x_13[15];
  assign wght_sign_x_13_16 = uSystolicPE_477_io_wght_sign_d;
  assign wght_abs_x_13_16 = uSystolicPE_477_io_wght_abs_d;
  assign uSystolicPE_477_io_enable_o = enable_o_x_13[16];
  assign uSystolicPE_477_io_clear_o = clear_o_x_13[16];
  assign ofm_x_13_15 = uSystolicPE_477_io_ofm_d;
  assign randW_x_15_14 = uSystolicPE_477_io_randW_d;
  assign uSystolicPE_478_io_mac_done = mac_done_x_15[14];
  assign uSystolicPE_478_io_enable_i = enable_i_x_15[14];
  assign uSystolicPE_478_io_clear_i = clear_i_x_15[14];
  assign ifm_sign_x_15_15 = uSystolicPE_478_io_ifm_sign_d;
  assign ifm_dff_x_15_15 = uSystolicPE_478_io_ifm_dff_d;
  assign uSystolicPE_478_io_enable_w = enable_w_x_14[15];
  assign uSystolicPE_478_io_clear_w = clear_w_x_14[15];
  assign wght_sign_x_14_16 = uSystolicPE_478_io_wght_sign_d;
  assign wght_abs_x_14_16 = uSystolicPE_478_io_wght_abs_d;
  assign uSystolicPE_478_io_enable_o = enable_o_x_14[16];
  assign uSystolicPE_478_io_clear_o = clear_o_x_14[16];
  assign ofm_x_14_15 = uSystolicPE_478_io_ofm_d;
  assign randW_x_15_15 = uSystolicPE_478_io_randW_d;
  assign uSystolicPE_479_io_mac_done = mac_done_x_15[15];
  assign uSystolicPE_479_io_enable_i = enable_i_x_15[15];
  assign uSystolicPE_479_io_clear_i = clear_i_x_15[15];
  assign ifm_sign_x_15_16 = uSystolicPE_479_io_ifm_sign_d;
  assign ifm_dff_x_15_16 = uSystolicPE_479_io_ifm_dff_d;
  assign uSystolicPE_479_io_enable_w = enable_w_x_15[15];
  assign uSystolicPE_479_io_clear_w = clear_w_x_15[15];
  assign wght_sign_x_15_16 = uSystolicPE_479_io_wght_sign_d;
  assign wght_abs_x_15_16 = uSystolicPE_479_io_wght_abs_d;
  assign uSystolicPE_479_io_enable_o = enable_o_x_15[16];
  assign uSystolicPE_479_io_clear_o = clear_o_x_15[16];
  assign ofm_x_15_15 = uSystolicPE_479_io_ofm_d;
  assign randW_x_15_16 = uSystolicPE_479_io_randW_d;

endmodule

//uSystolicPE_239 replaced by uSystolicPE

//uSystolicPE_238 replaced by uSystolicPE

//uSystolicPE_237 replaced by uSystolicPE

//uSystolicPE_236 replaced by uSystolicPE

//uSystolicPE_235 replaced by uSystolicPE

//uSystolicPE_234 replaced by uSystolicPE

//uSystolicPE_233 replaced by uSystolicPE

//uSystolicPE_232 replaced by uSystolicPE

//uSystolicPE_231 replaced by uSystolicPE

//uSystolicPE_230 replaced by uSystolicPE

//uSystolicPE_229 replaced by uSystolicPE

//uSystolicPE_228 replaced by uSystolicPE

//uSystolicPE_227 replaced by uSystolicPE

//uSystolicPE_226 replaced by uSystolicPE

//uSystolicPE_225 replaced by uSystolicPE

//uSystolicPEBorder_15 replaced by uSystolicPEBorder

//uSystolicPE_224 replaced by uSystolicPE

//uSystolicPE_223 replaced by uSystolicPE

//uSystolicPE_222 replaced by uSystolicPE

//uSystolicPE_221 replaced by uSystolicPE

//uSystolicPE_220 replaced by uSystolicPE

//uSystolicPE_219 replaced by uSystolicPE

//uSystolicPE_218 replaced by uSystolicPE

//uSystolicPE_217 replaced by uSystolicPE

//uSystolicPE_216 replaced by uSystolicPE

//uSystolicPE_215 replaced by uSystolicPE

//uSystolicPE_214 replaced by uSystolicPE

//uSystolicPE_213 replaced by uSystolicPE

//uSystolicPE_212 replaced by uSystolicPE

//uSystolicPE_211 replaced by uSystolicPE

//uSystolicPE_210 replaced by uSystolicPE

//uSystolicPEBorder_14 replaced by uSystolicPEBorder

//uSystolicPE_209 replaced by uSystolicPE

//uSystolicPE_208 replaced by uSystolicPE

//uSystolicPE_207 replaced by uSystolicPE

//uSystolicPE_206 replaced by uSystolicPE

//uSystolicPE_205 replaced by uSystolicPE

//uSystolicPE_204 replaced by uSystolicPE

//uSystolicPE_203 replaced by uSystolicPE

//uSystolicPE_202 replaced by uSystolicPE

//uSystolicPE_201 replaced by uSystolicPE

//uSystolicPE_200 replaced by uSystolicPE

//uSystolicPE_199 replaced by uSystolicPE

//uSystolicPE_198 replaced by uSystolicPE

//uSystolicPE_197 replaced by uSystolicPE

//uSystolicPE_196 replaced by uSystolicPE

//uSystolicPE_195 replaced by uSystolicPE

//uSystolicPEBorder_13 replaced by uSystolicPEBorder

//uSystolicPE_194 replaced by uSystolicPE

//uSystolicPE_193 replaced by uSystolicPE

//uSystolicPE_192 replaced by uSystolicPE

//uSystolicPE_191 replaced by uSystolicPE

//uSystolicPE_190 replaced by uSystolicPE

//uSystolicPE_189 replaced by uSystolicPE

//uSystolicPE_188 replaced by uSystolicPE

//uSystolicPE_187 replaced by uSystolicPE

//uSystolicPE_186 replaced by uSystolicPE

//uSystolicPE_185 replaced by uSystolicPE

//uSystolicPE_184 replaced by uSystolicPE

//uSystolicPE_183 replaced by uSystolicPE

//uSystolicPE_182 replaced by uSystolicPE

//uSystolicPE_181 replaced by uSystolicPE

//uSystolicPE_180 replaced by uSystolicPE

//uSystolicPEBorder_12 replaced by uSystolicPEBorder

//uSystolicPE_179 replaced by uSystolicPE

//uSystolicPE_178 replaced by uSystolicPE

//uSystolicPE_177 replaced by uSystolicPE

//uSystolicPE_176 replaced by uSystolicPE

//uSystolicPE_175 replaced by uSystolicPE

//uSystolicPE_174 replaced by uSystolicPE

//uSystolicPE_173 replaced by uSystolicPE

//uSystolicPE_172 replaced by uSystolicPE

//uSystolicPE_171 replaced by uSystolicPE

//uSystolicPE_170 replaced by uSystolicPE

//uSystolicPE_169 replaced by uSystolicPE

//uSystolicPE_168 replaced by uSystolicPE

//uSystolicPE_167 replaced by uSystolicPE

//uSystolicPE_166 replaced by uSystolicPE

//uSystolicPE_165 replaced by uSystolicPE

//uSystolicPEBorder_11 replaced by uSystolicPEBorder

//uSystolicPE_164 replaced by uSystolicPE

//uSystolicPE_163 replaced by uSystolicPE

//uSystolicPE_162 replaced by uSystolicPE

//uSystolicPE_161 replaced by uSystolicPE

//uSystolicPE_160 replaced by uSystolicPE

//uSystolicPE_159 replaced by uSystolicPE

//uSystolicPE_158 replaced by uSystolicPE

//uSystolicPE_157 replaced by uSystolicPE

//uSystolicPE_156 replaced by uSystolicPE

//uSystolicPE_155 replaced by uSystolicPE

//uSystolicPE_154 replaced by uSystolicPE

//uSystolicPE_153 replaced by uSystolicPE

//uSystolicPE_152 replaced by uSystolicPE

//uSystolicPE_151 replaced by uSystolicPE

//uSystolicPE_150 replaced by uSystolicPE

//uSystolicPEBorder_10 replaced by uSystolicPEBorder

//uSystolicPE_149 replaced by uSystolicPE

//uSystolicPE_148 replaced by uSystolicPE

//uSystolicPE_147 replaced by uSystolicPE

//uSystolicPE_146 replaced by uSystolicPE

//uSystolicPE_145 replaced by uSystolicPE

//uSystolicPE_144 replaced by uSystolicPE

//uSystolicPE_143 replaced by uSystolicPE

//uSystolicPE_142 replaced by uSystolicPE

//uSystolicPE_141 replaced by uSystolicPE

//uSystolicPE_140 replaced by uSystolicPE

//uSystolicPE_139 replaced by uSystolicPE

//uSystolicPE_138 replaced by uSystolicPE

//uSystolicPE_137 replaced by uSystolicPE

//uSystolicPE_136 replaced by uSystolicPE

//uSystolicPE_135 replaced by uSystolicPE

//uSystolicPEBorder_9 replaced by uSystolicPEBorder

//uSystolicPE_134 replaced by uSystolicPE

//uSystolicPE_133 replaced by uSystolicPE

//uSystolicPE_132 replaced by uSystolicPE

//uSystolicPE_131 replaced by uSystolicPE

//uSystolicPE_130 replaced by uSystolicPE

//uSystolicPE_129 replaced by uSystolicPE

//uSystolicPE_128 replaced by uSystolicPE

//uSystolicPE_127 replaced by uSystolicPE

//uSystolicPE_126 replaced by uSystolicPE

//uSystolicPE_125 replaced by uSystolicPE

//uSystolicPE_124 replaced by uSystolicPE

//uSystolicPE_123 replaced by uSystolicPE

//uSystolicPE_122 replaced by uSystolicPE

//uSystolicPE_121 replaced by uSystolicPE

//uSystolicPE_120 replaced by uSystolicPE

//uSystolicPEBorder_8 replaced by uSystolicPEBorder

//uSystolicPE_119 replaced by uSystolicPE

//uSystolicPE_118 replaced by uSystolicPE

//uSystolicPE_117 replaced by uSystolicPE

//uSystolicPE_116 replaced by uSystolicPE

//uSystolicPE_115 replaced by uSystolicPE

//uSystolicPE_114 replaced by uSystolicPE

//uSystolicPE_113 replaced by uSystolicPE

//uSystolicPE_112 replaced by uSystolicPE

//uSystolicPE_111 replaced by uSystolicPE

//uSystolicPE_110 replaced by uSystolicPE

//uSystolicPE_109 replaced by uSystolicPE

//uSystolicPE_108 replaced by uSystolicPE

//uSystolicPE_107 replaced by uSystolicPE

//uSystolicPE_106 replaced by uSystolicPE

//uSystolicPE_105 replaced by uSystolicPE

//uSystolicPEBorder_7 replaced by uSystolicPEBorder

//uSystolicPE_104 replaced by uSystolicPE

//uSystolicPE_103 replaced by uSystolicPE

//uSystolicPE_102 replaced by uSystolicPE

//uSystolicPE_101 replaced by uSystolicPE

//uSystolicPE_100 replaced by uSystolicPE

//uSystolicPE_99 replaced by uSystolicPE

//uSystolicPE_98 replaced by uSystolicPE

//uSystolicPE_97 replaced by uSystolicPE

//uSystolicPE_96 replaced by uSystolicPE

//uSystolicPE_95 replaced by uSystolicPE

//uSystolicPE_94 replaced by uSystolicPE

//uSystolicPE_93 replaced by uSystolicPE

//uSystolicPE_92 replaced by uSystolicPE

//uSystolicPE_91 replaced by uSystolicPE

//uSystolicPE_90 replaced by uSystolicPE

//uSystolicPEBorder_6 replaced by uSystolicPEBorder

//uSystolicPE_89 replaced by uSystolicPE

//uSystolicPE_88 replaced by uSystolicPE

//uSystolicPE_87 replaced by uSystolicPE

//uSystolicPE_86 replaced by uSystolicPE

//uSystolicPE_85 replaced by uSystolicPE

//uSystolicPE_84 replaced by uSystolicPE

//uSystolicPE_83 replaced by uSystolicPE

//uSystolicPE_82 replaced by uSystolicPE

//uSystolicPE_81 replaced by uSystolicPE

//uSystolicPE_80 replaced by uSystolicPE

//uSystolicPE_79 replaced by uSystolicPE

//uSystolicPE_78 replaced by uSystolicPE

//uSystolicPE_77 replaced by uSystolicPE

//uSystolicPE_76 replaced by uSystolicPE

//uSystolicPE_75 replaced by uSystolicPE

//uSystolicPEBorder_5 replaced by uSystolicPEBorder

//uSystolicPE_74 replaced by uSystolicPE

//uSystolicPE_73 replaced by uSystolicPE

//uSystolicPE_72 replaced by uSystolicPE

//uSystolicPE_71 replaced by uSystolicPE

//uSystolicPE_70 replaced by uSystolicPE

//uSystolicPE_69 replaced by uSystolicPE

//uSystolicPE_68 replaced by uSystolicPE

//uSystolicPE_67 replaced by uSystolicPE

//uSystolicPE_66 replaced by uSystolicPE

//uSystolicPE_65 replaced by uSystolicPE

//uSystolicPE_64 replaced by uSystolicPE

//uSystolicPE_63 replaced by uSystolicPE

//uSystolicPE_62 replaced by uSystolicPE

//uSystolicPE_61 replaced by uSystolicPE

//uSystolicPE_60 replaced by uSystolicPE

//uSystolicPEBorder_4 replaced by uSystolicPEBorder

//uSystolicPE_59 replaced by uSystolicPE

//uSystolicPE_58 replaced by uSystolicPE

//uSystolicPE_57 replaced by uSystolicPE

//uSystolicPE_56 replaced by uSystolicPE

//uSystolicPE_55 replaced by uSystolicPE

//uSystolicPE_54 replaced by uSystolicPE

//uSystolicPE_53 replaced by uSystolicPE

//uSystolicPE_52 replaced by uSystolicPE

//uSystolicPE_51 replaced by uSystolicPE

//uSystolicPE_50 replaced by uSystolicPE

//uSystolicPE_49 replaced by uSystolicPE

//uSystolicPE_48 replaced by uSystolicPE

//uSystolicPE_47 replaced by uSystolicPE

//uSystolicPE_46 replaced by uSystolicPE

//uSystolicPE_45 replaced by uSystolicPE

//uSystolicPEBorder_3 replaced by uSystolicPEBorder

//uSystolicPE_44 replaced by uSystolicPE

//uSystolicPE_43 replaced by uSystolicPE

//uSystolicPE_42 replaced by uSystolicPE

//uSystolicPE_41 replaced by uSystolicPE

//uSystolicPE_40 replaced by uSystolicPE

//uSystolicPE_39 replaced by uSystolicPE

//uSystolicPE_38 replaced by uSystolicPE

//uSystolicPE_37 replaced by uSystolicPE

//uSystolicPE_36 replaced by uSystolicPE

//uSystolicPE_35 replaced by uSystolicPE

//uSystolicPE_34 replaced by uSystolicPE

//uSystolicPE_33 replaced by uSystolicPE

//uSystolicPE_32 replaced by uSystolicPE

//uSystolicPE_31 replaced by uSystolicPE

//uSystolicPE_30 replaced by uSystolicPE

//uSystolicPEBorder_2 replaced by uSystolicPEBorder

//uSystolicPE_29 replaced by uSystolicPE

//uSystolicPE_28 replaced by uSystolicPE

//uSystolicPE_27 replaced by uSystolicPE

//uSystolicPE_26 replaced by uSystolicPE

//uSystolicPE_25 replaced by uSystolicPE

//uSystolicPE_24 replaced by uSystolicPE

//uSystolicPE_23 replaced by uSystolicPE

//uSystolicPE_22 replaced by uSystolicPE

//uSystolicPE_21 replaced by uSystolicPE

//uSystolicPE_20 replaced by uSystolicPE

//uSystolicPE_19 replaced by uSystolicPE

//uSystolicPE_18 replaced by uSystolicPE

//uSystolicPE_17 replaced by uSystolicPE

//uSystolicPE_16 replaced by uSystolicPE

//uSystolicPE_15 replaced by uSystolicPE

//uSystolicPEBorder_1 replaced by uSystolicPEBorder

//uSystolicPE_14 replaced by uSystolicPE

//uSystolicPE_13 replaced by uSystolicPE

//uSystolicPE_12 replaced by uSystolicPE

//uSystolicPE_11 replaced by uSystolicPE

//uSystolicPE_10 replaced by uSystolicPE

//uSystolicPE_9 replaced by uSystolicPE

//uSystolicPE_8 replaced by uSystolicPE

//uSystolicPE_7 replaced by uSystolicPE

//uSystolicPE_6 replaced by uSystolicPE

//uSystolicPE_5 replaced by uSystolicPE

//uSystolicPE_4 replaced by uSystolicPE

//uSystolicPE_3 replaced by uSystolicPE

//uSystolicPE_2 replaced by uSystolicPE

//uSystolicPE_1 replaced by uSystolicPE

module uSystolicPE (
  input  wire          io_mac_done,
  input  wire          io_enable_i,
  input  wire          io_clear_i,
  input  wire          io_enable_w,
  input  wire          io_clear_w,
  input  wire          io_enable_o,
  input  wire          io_clear_o,
  input  wire          io_ifm_sign,
  input  wire          io_ifm_dff,
  input  wire          io_wght_sign,
  input  wire [14:0]   io_randW,
  input  wire [14:0]   io_wght_abs,
  input  wire [31:0]   io_ofm,
  output wire          io_mac_done_d,
  output wire          io_enable_i_d,
  output wire          io_clear_i_d,
  output wire          io_enable_w_d,
  output wire          io_clear_w_d,
  output wire          io_enable_o_d,
  output wire          io_clear_o_d,
  output wire          io_ifm_sign_d,
  output wire          io_ifm_dff_d,
  output wire          io_wght_sign_d,
  output wire [14:0]   io_randW_d,
  output wire [14:0]   io_wght_abs_d,
  output wire [31:0]   io_ofm_d,
  input  wire          clk,
  input  wire          reset
);

  wire                ireg_inner_io_o_data_sign;
  wire                ireg_inner_io_o_data_dff;
  wire       [14:0]   wreg_inner_io_output_abs;
  wire                wreg_inner_io_output_sign;
  wire       [14:0]   umul_inner_io_o_randw;
  wire                umul_inner_io_o_bit;
  wire       [31:0]   acc_io_sum_output;

  ireg_239 ireg_inner (
    .io_enable      (io_enable_i              ), //i
    .io_clear       (io_clear_i               ), //i
    .io_i_data_sign (io_ifm_sign              ), //i
    .io_i_data_dff  (io_ifm_dff               ), //i
    .io_o_data_sign (ireg_inner_io_o_data_sign), //o
    .io_o_data_dff  (ireg_inner_io_o_data_dff ), //o
    .clk            (clk                      ), //i
    .reset          (reset                    )  //i
  );
  wreg_255 wreg_inner (
    .io_enable      (io_enable_w                   ), //i
    .io_clear       (io_clear_w                    ), //i
    .io_input_abs   (io_wght_abs[14:0]             ), //i
    .io_input_sign  (io_wght_sign                  ), //i
    .io_output_abs  (wreg_inner_io_output_abs[14:0]), //o
    .io_output_sign (wreg_inner_io_output_sign     ), //o
    .clk            (clk                           ), //i
    .reset          (reset                         )  //i
  );
  umul_239 umul_inner (
    .io_i_bit_i  (io_ifm_dff_d               ), //i
    .io_i_data_w (io_wght_abs_d[14:0]        ), //i
    .io_i_randw  (io_randW[14:0]             ), //i
    .io_o_randw  (umul_inner_io_o_randw[14:0]), //o
    .io_o_bit    (umul_inner_io_o_bit        )  //o
  );
  accumulate_255 acc (
    .io_enable          (io_enable_o            ), //i
    .io_clear           (io_clear_o             ), //i
    .io_mac_done        (io_mac_done_d          ), //i
    .io_sign_activation (io_ifm_sign_d          ), //i
    .io_sign_weight     (io_wght_sign_d         ), //i
    .io_sum_input       (io_ofm[31:0]           ), //i
    .io_sum_output      (acc_io_sum_output[31:0]), //o
    .io_prod_bit        (umul_inner_io_o_bit    ), //i
    .clk                (clk                    ), //i
    .reset              (reset                  )  //i
  );
  assign io_ifm_sign_d = ireg_inner_io_o_data_sign;
  assign io_ifm_dff_d = ireg_inner_io_o_data_dff;
  assign io_wght_sign_d = wreg_inner_io_output_sign;
  assign io_wght_abs_d = wreg_inner_io_output_abs;
  assign io_randW_d = umul_inner_io_o_randw;
  assign io_ofm_d = acc_io_sum_output;
  assign io_enable_i_d = io_enable_i;
  assign io_enable_w_d = io_enable_w;
  assign io_enable_o_d = io_enable_o;
  assign io_clear_i_d = io_clear_i;
  assign io_clear_w_d = io_clear_w;
  assign io_clear_o_d = io_clear_o;
  assign io_mac_done_d = io_mac_done;

endmodule

module uSystolicPEBorder (
  input  wire          io_mac_done,
  input  wire          io_enable_i,
  input  wire          io_clear_i,
  input  wire          io_enable_w,
  input  wire          io_clear_w,
  input  wire          io_enable_o,
  input  wire          io_clear_o,
  input  wire [15:0]   io_ifm,
  input  wire          io_wght_sign,
  input  wire [14:0]   io_wght_abs,
  input  wire [31:0]   io_ofm,
  output wire          io_mac_done_d,
  output wire          io_enable_i_d,
  output wire          io_clear_i_d,
  output wire          io_enable_w_d,
  output wire          io_clear_w_d,
  output wire          io_enable_o_d,
  output wire          io_clear_o_d,
  output wire          io_ifm_sign_d,
  output wire          io_ifm_dff_d,
  output wire          io_wght_sign_d,
  output wire [14:0]   io_randW_d,
  output wire [14:0]   io_wght_abs_d,
  output wire [31:0]   io_ofm_d,
  input  wire          clk,
  input  wire          reset
);

  wire                ireg_border_io_output_sign;
  wire       [14:0]   ireg_border_io_output_abs;
  wire       [14:0]   wreg_border_io_output_abs;
  wire                wreg_border_io_output_sign;
  wire       [14:0]   umul_border_io_randW;
  wire                umul_border_io_o_bit;
  wire                umul_border_io_i_bit_d;
  wire       [31:0]   acc_io_sum_output;

  uregBorder_15 ireg_border (
    .io_enable      (io_enable_i                    ), //i
    .io_clear       (io_clear_i                     ), //i
    .io_input       (io_ifm[15:0]                   ), //i
    .io_output_sign (ireg_border_io_output_sign     ), //o
    .io_output_abs  (ireg_border_io_output_abs[14:0]), //o
    .clk            (clk                            ), //i
    .reset          (reset                          )  //i
  );
  wreg_255 wreg_border (
    .io_enable      (io_enable_w                    ), //i
    .io_clear       (io_clear_w                     ), //i
    .io_input_abs   (io_wght_abs[14:0]              ), //i
    .io_input_sign  (io_wght_sign                   ), //i
    .io_output_abs  (wreg_border_io_output_abs[14:0]), //o
    .io_output_sign (wreg_border_io_output_sign     ), //o
    .clk            (clk                            ), //i
    .reset          (reset                          )  //i
  );
  umulBorder_15 umul_border (
    .io_clear    (io_clear_i_d                   ), //i
    .io_init     (io_enable_i_d                  ), //i
    .io_i_data_i (ireg_border_io_output_abs[14:0]), //i
    .io_i_data_w (io_wght_abs_d[14:0]            ), //i
    .io_randW    (umul_border_io_randW[14:0]     ), //o
    .io_o_bit    (umul_border_io_o_bit           ), //o
    .io_i_bit_d  (umul_border_io_i_bit_d         ), //o
    .clk         (clk                            ), //i
    .reset       (reset                          )  //i
  );
  accumulate_255 acc (
    .io_enable          (io_enable_o            ), //i
    .io_clear           (io_clear_o             ), //i
    .io_mac_done        (io_mac_done_d          ), //i
    .io_sign_activation (io_ifm_sign_d          ), //i
    .io_sign_weight     (io_wght_sign_d         ), //i
    .io_sum_input       (io_ofm[31:0]           ), //i
    .io_sum_output      (acc_io_sum_output[31:0]), //o
    .io_prod_bit        (umul_border_io_o_bit   ), //i
    .clk                (clk                    ), //i
    .reset              (reset                  )  //i
  );
  assign io_ifm_sign_d = ireg_border_io_output_sign;
  assign io_wght_sign_d = wreg_border_io_output_sign;
  assign io_wght_abs_d = wreg_border_io_output_abs;
  assign io_randW_d = umul_border_io_randW;
  assign io_ifm_dff_d = umul_border_io_i_bit_d;
  assign io_ofm_d = acc_io_sum_output;
  assign io_enable_i_d = io_enable_i;
  assign io_enable_w_d = io_enable_w;
  assign io_enable_o_d = io_enable_o;
  assign io_clear_i_d = io_clear_i;
  assign io_clear_w_d = io_clear_w;
  assign io_clear_o_d = io_clear_o;
  assign io_mac_done_d = io_mac_done;

endmodule

//accumulate replaced by accumulate_255

//umul replaced by umul_239

//wreg replaced by wreg_255

//ireg replaced by ireg_239

//accumulate_1 replaced by accumulate_255

//umul_1 replaced by umul_239

//wreg_1 replaced by wreg_255

//ireg_1 replaced by ireg_239

//accumulate_2 replaced by accumulate_255

//umul_2 replaced by umul_239

//wreg_2 replaced by wreg_255

//ireg_2 replaced by ireg_239

//accumulate_3 replaced by accumulate_255

//umul_3 replaced by umul_239

//wreg_3 replaced by wreg_255

//ireg_3 replaced by ireg_239

//accumulate_4 replaced by accumulate_255

//umul_4 replaced by umul_239

//wreg_4 replaced by wreg_255

//ireg_4 replaced by ireg_239

//accumulate_5 replaced by accumulate_255

//umul_5 replaced by umul_239

//wreg_5 replaced by wreg_255

//ireg_5 replaced by ireg_239

//accumulate_6 replaced by accumulate_255

//umul_6 replaced by umul_239

//wreg_6 replaced by wreg_255

//ireg_6 replaced by ireg_239

//accumulate_7 replaced by accumulate_255

//umul_7 replaced by umul_239

//wreg_7 replaced by wreg_255

//ireg_7 replaced by ireg_239

//accumulate_8 replaced by accumulate_255

//umul_8 replaced by umul_239

//wreg_8 replaced by wreg_255

//ireg_8 replaced by ireg_239

//accumulate_9 replaced by accumulate_255

//umul_9 replaced by umul_239

//wreg_9 replaced by wreg_255

//ireg_9 replaced by ireg_239

//accumulate_10 replaced by accumulate_255

//umul_10 replaced by umul_239

//wreg_10 replaced by wreg_255

//ireg_10 replaced by ireg_239

//accumulate_11 replaced by accumulate_255

//umul_11 replaced by umul_239

//wreg_11 replaced by wreg_255

//ireg_11 replaced by ireg_239

//accumulate_12 replaced by accumulate_255

//umul_12 replaced by umul_239

//wreg_12 replaced by wreg_255

//ireg_12 replaced by ireg_239

//accumulate_13 replaced by accumulate_255

//umul_13 replaced by umul_239

//wreg_13 replaced by wreg_255

//ireg_13 replaced by ireg_239

//accumulate_14 replaced by accumulate_255

//umul_14 replaced by umul_239

//wreg_14 replaced by wreg_255

//ireg_14 replaced by ireg_239

//accumulate_15 replaced by accumulate_255

//umulBorder replaced by umulBorder_15

//wreg_15 replaced by wreg_255

//uregBorder replaced by uregBorder_15

//accumulate_16 replaced by accumulate_255

//umul_15 replaced by umul_239

//wreg_16 replaced by wreg_255

//ireg_15 replaced by ireg_239

//accumulate_17 replaced by accumulate_255

//umul_16 replaced by umul_239

//wreg_17 replaced by wreg_255

//ireg_16 replaced by ireg_239

//accumulate_18 replaced by accumulate_255

//umul_17 replaced by umul_239

//wreg_18 replaced by wreg_255

//ireg_17 replaced by ireg_239

//accumulate_19 replaced by accumulate_255

//umul_18 replaced by umul_239

//wreg_19 replaced by wreg_255

//ireg_18 replaced by ireg_239

//accumulate_20 replaced by accumulate_255

//umul_19 replaced by umul_239

//wreg_20 replaced by wreg_255

//ireg_19 replaced by ireg_239

//accumulate_21 replaced by accumulate_255

//umul_20 replaced by umul_239

//wreg_21 replaced by wreg_255

//ireg_20 replaced by ireg_239

//accumulate_22 replaced by accumulate_255

//umul_21 replaced by umul_239

//wreg_22 replaced by wreg_255

//ireg_21 replaced by ireg_239

//accumulate_23 replaced by accumulate_255

//umul_22 replaced by umul_239

//wreg_23 replaced by wreg_255

//ireg_22 replaced by ireg_239

//accumulate_24 replaced by accumulate_255

//umul_23 replaced by umul_239

//wreg_24 replaced by wreg_255

//ireg_23 replaced by ireg_239

//accumulate_25 replaced by accumulate_255

//umul_24 replaced by umul_239

//wreg_25 replaced by wreg_255

//ireg_24 replaced by ireg_239

//accumulate_26 replaced by accumulate_255

//umul_25 replaced by umul_239

//wreg_26 replaced by wreg_255

//ireg_25 replaced by ireg_239

//accumulate_27 replaced by accumulate_255

//umul_26 replaced by umul_239

//wreg_27 replaced by wreg_255

//ireg_26 replaced by ireg_239

//accumulate_28 replaced by accumulate_255

//umul_27 replaced by umul_239

//wreg_28 replaced by wreg_255

//ireg_27 replaced by ireg_239

//accumulate_29 replaced by accumulate_255

//umul_28 replaced by umul_239

//wreg_29 replaced by wreg_255

//ireg_28 replaced by ireg_239

//accumulate_30 replaced by accumulate_255

//umul_29 replaced by umul_239

//wreg_30 replaced by wreg_255

//ireg_29 replaced by ireg_239

//accumulate_31 replaced by accumulate_255

//umulBorder_1 replaced by umulBorder_15

//wreg_31 replaced by wreg_255

//uregBorder_1 replaced by uregBorder_15

//accumulate_32 replaced by accumulate_255

//umul_30 replaced by umul_239

//wreg_32 replaced by wreg_255

//ireg_30 replaced by ireg_239

//accumulate_33 replaced by accumulate_255

//umul_31 replaced by umul_239

//wreg_33 replaced by wreg_255

//ireg_31 replaced by ireg_239

//accumulate_34 replaced by accumulate_255

//umul_32 replaced by umul_239

//wreg_34 replaced by wreg_255

//ireg_32 replaced by ireg_239

//accumulate_35 replaced by accumulate_255

//umul_33 replaced by umul_239

//wreg_35 replaced by wreg_255

//ireg_33 replaced by ireg_239

//accumulate_36 replaced by accumulate_255

//umul_34 replaced by umul_239

//wreg_36 replaced by wreg_255

//ireg_34 replaced by ireg_239

//accumulate_37 replaced by accumulate_255

//umul_35 replaced by umul_239

//wreg_37 replaced by wreg_255

//ireg_35 replaced by ireg_239

//accumulate_38 replaced by accumulate_255

//umul_36 replaced by umul_239

//wreg_38 replaced by wreg_255

//ireg_36 replaced by ireg_239

//accumulate_39 replaced by accumulate_255

//umul_37 replaced by umul_239

//wreg_39 replaced by wreg_255

//ireg_37 replaced by ireg_239

//accumulate_40 replaced by accumulate_255

//umul_38 replaced by umul_239

//wreg_40 replaced by wreg_255

//ireg_38 replaced by ireg_239

//accumulate_41 replaced by accumulate_255

//umul_39 replaced by umul_239

//wreg_41 replaced by wreg_255

//ireg_39 replaced by ireg_239

//accumulate_42 replaced by accumulate_255

//umul_40 replaced by umul_239

//wreg_42 replaced by wreg_255

//ireg_40 replaced by ireg_239

//accumulate_43 replaced by accumulate_255

//umul_41 replaced by umul_239

//wreg_43 replaced by wreg_255

//ireg_41 replaced by ireg_239

//accumulate_44 replaced by accumulate_255

//umul_42 replaced by umul_239

//wreg_44 replaced by wreg_255

//ireg_42 replaced by ireg_239

//accumulate_45 replaced by accumulate_255

//umul_43 replaced by umul_239

//wreg_45 replaced by wreg_255

//ireg_43 replaced by ireg_239

//accumulate_46 replaced by accumulate_255

//umul_44 replaced by umul_239

//wreg_46 replaced by wreg_255

//ireg_44 replaced by ireg_239

//accumulate_47 replaced by accumulate_255

//umulBorder_2 replaced by umulBorder_15

//wreg_47 replaced by wreg_255

//uregBorder_2 replaced by uregBorder_15

//accumulate_48 replaced by accumulate_255

//umul_45 replaced by umul_239

//wreg_48 replaced by wreg_255

//ireg_45 replaced by ireg_239

//accumulate_49 replaced by accumulate_255

//umul_46 replaced by umul_239

//wreg_49 replaced by wreg_255

//ireg_46 replaced by ireg_239

//accumulate_50 replaced by accumulate_255

//umul_47 replaced by umul_239

//wreg_50 replaced by wreg_255

//ireg_47 replaced by ireg_239

//accumulate_51 replaced by accumulate_255

//umul_48 replaced by umul_239

//wreg_51 replaced by wreg_255

//ireg_48 replaced by ireg_239

//accumulate_52 replaced by accumulate_255

//umul_49 replaced by umul_239

//wreg_52 replaced by wreg_255

//ireg_49 replaced by ireg_239

//accumulate_53 replaced by accumulate_255

//umul_50 replaced by umul_239

//wreg_53 replaced by wreg_255

//ireg_50 replaced by ireg_239

//accumulate_54 replaced by accumulate_255

//umul_51 replaced by umul_239

//wreg_54 replaced by wreg_255

//ireg_51 replaced by ireg_239

//accumulate_55 replaced by accumulate_255

//umul_52 replaced by umul_239

//wreg_55 replaced by wreg_255

//ireg_52 replaced by ireg_239

//accumulate_56 replaced by accumulate_255

//umul_53 replaced by umul_239

//wreg_56 replaced by wreg_255

//ireg_53 replaced by ireg_239

//accumulate_57 replaced by accumulate_255

//umul_54 replaced by umul_239

//wreg_57 replaced by wreg_255

//ireg_54 replaced by ireg_239

//accumulate_58 replaced by accumulate_255

//umul_55 replaced by umul_239

//wreg_58 replaced by wreg_255

//ireg_55 replaced by ireg_239

//accumulate_59 replaced by accumulate_255

//umul_56 replaced by umul_239

//wreg_59 replaced by wreg_255

//ireg_56 replaced by ireg_239

//accumulate_60 replaced by accumulate_255

//umul_57 replaced by umul_239

//wreg_60 replaced by wreg_255

//ireg_57 replaced by ireg_239

//accumulate_61 replaced by accumulate_255

//umul_58 replaced by umul_239

//wreg_61 replaced by wreg_255

//ireg_58 replaced by ireg_239

//accumulate_62 replaced by accumulate_255

//umul_59 replaced by umul_239

//wreg_62 replaced by wreg_255

//ireg_59 replaced by ireg_239

//accumulate_63 replaced by accumulate_255

//umulBorder_3 replaced by umulBorder_15

//wreg_63 replaced by wreg_255

//uregBorder_3 replaced by uregBorder_15

//accumulate_64 replaced by accumulate_255

//umul_60 replaced by umul_239

//wreg_64 replaced by wreg_255

//ireg_60 replaced by ireg_239

//accumulate_65 replaced by accumulate_255

//umul_61 replaced by umul_239

//wreg_65 replaced by wreg_255

//ireg_61 replaced by ireg_239

//accumulate_66 replaced by accumulate_255

//umul_62 replaced by umul_239

//wreg_66 replaced by wreg_255

//ireg_62 replaced by ireg_239

//accumulate_67 replaced by accumulate_255

//umul_63 replaced by umul_239

//wreg_67 replaced by wreg_255

//ireg_63 replaced by ireg_239

//accumulate_68 replaced by accumulate_255

//umul_64 replaced by umul_239

//wreg_68 replaced by wreg_255

//ireg_64 replaced by ireg_239

//accumulate_69 replaced by accumulate_255

//umul_65 replaced by umul_239

//wreg_69 replaced by wreg_255

//ireg_65 replaced by ireg_239

//accumulate_70 replaced by accumulate_255

//umul_66 replaced by umul_239

//wreg_70 replaced by wreg_255

//ireg_66 replaced by ireg_239

//accumulate_71 replaced by accumulate_255

//umul_67 replaced by umul_239

//wreg_71 replaced by wreg_255

//ireg_67 replaced by ireg_239

//accumulate_72 replaced by accumulate_255

//umul_68 replaced by umul_239

//wreg_72 replaced by wreg_255

//ireg_68 replaced by ireg_239

//accumulate_73 replaced by accumulate_255

//umul_69 replaced by umul_239

//wreg_73 replaced by wreg_255

//ireg_69 replaced by ireg_239

//accumulate_74 replaced by accumulate_255

//umul_70 replaced by umul_239

//wreg_74 replaced by wreg_255

//ireg_70 replaced by ireg_239

//accumulate_75 replaced by accumulate_255

//umul_71 replaced by umul_239

//wreg_75 replaced by wreg_255

//ireg_71 replaced by ireg_239

//accumulate_76 replaced by accumulate_255

//umul_72 replaced by umul_239

//wreg_76 replaced by wreg_255

//ireg_72 replaced by ireg_239

//accumulate_77 replaced by accumulate_255

//umul_73 replaced by umul_239

//wreg_77 replaced by wreg_255

//ireg_73 replaced by ireg_239

//accumulate_78 replaced by accumulate_255

//umul_74 replaced by umul_239

//wreg_78 replaced by wreg_255

//ireg_74 replaced by ireg_239

//accumulate_79 replaced by accumulate_255

//umulBorder_4 replaced by umulBorder_15

//wreg_79 replaced by wreg_255

//uregBorder_4 replaced by uregBorder_15

//accumulate_80 replaced by accumulate_255

//umul_75 replaced by umul_239

//wreg_80 replaced by wreg_255

//ireg_75 replaced by ireg_239

//accumulate_81 replaced by accumulate_255

//umul_76 replaced by umul_239

//wreg_81 replaced by wreg_255

//ireg_76 replaced by ireg_239

//accumulate_82 replaced by accumulate_255

//umul_77 replaced by umul_239

//wreg_82 replaced by wreg_255

//ireg_77 replaced by ireg_239

//accumulate_83 replaced by accumulate_255

//umul_78 replaced by umul_239

//wreg_83 replaced by wreg_255

//ireg_78 replaced by ireg_239

//accumulate_84 replaced by accumulate_255

//umul_79 replaced by umul_239

//wreg_84 replaced by wreg_255

//ireg_79 replaced by ireg_239

//accumulate_85 replaced by accumulate_255

//umul_80 replaced by umul_239

//wreg_85 replaced by wreg_255

//ireg_80 replaced by ireg_239

//accumulate_86 replaced by accumulate_255

//umul_81 replaced by umul_239

//wreg_86 replaced by wreg_255

//ireg_81 replaced by ireg_239

//accumulate_87 replaced by accumulate_255

//umul_82 replaced by umul_239

//wreg_87 replaced by wreg_255

//ireg_82 replaced by ireg_239

//accumulate_88 replaced by accumulate_255

//umul_83 replaced by umul_239

//wreg_88 replaced by wreg_255

//ireg_83 replaced by ireg_239

//accumulate_89 replaced by accumulate_255

//umul_84 replaced by umul_239

//wreg_89 replaced by wreg_255

//ireg_84 replaced by ireg_239

//accumulate_90 replaced by accumulate_255

//umul_85 replaced by umul_239

//wreg_90 replaced by wreg_255

//ireg_85 replaced by ireg_239

//accumulate_91 replaced by accumulate_255

//umul_86 replaced by umul_239

//wreg_91 replaced by wreg_255

//ireg_86 replaced by ireg_239

//accumulate_92 replaced by accumulate_255

//umul_87 replaced by umul_239

//wreg_92 replaced by wreg_255

//ireg_87 replaced by ireg_239

//accumulate_93 replaced by accumulate_255

//umul_88 replaced by umul_239

//wreg_93 replaced by wreg_255

//ireg_88 replaced by ireg_239

//accumulate_94 replaced by accumulate_255

//umul_89 replaced by umul_239

//wreg_94 replaced by wreg_255

//ireg_89 replaced by ireg_239

//accumulate_95 replaced by accumulate_255

//umulBorder_5 replaced by umulBorder_15

//wreg_95 replaced by wreg_255

//uregBorder_5 replaced by uregBorder_15

//accumulate_96 replaced by accumulate_255

//umul_90 replaced by umul_239

//wreg_96 replaced by wreg_255

//ireg_90 replaced by ireg_239

//accumulate_97 replaced by accumulate_255

//umul_91 replaced by umul_239

//wreg_97 replaced by wreg_255

//ireg_91 replaced by ireg_239

//accumulate_98 replaced by accumulate_255

//umul_92 replaced by umul_239

//wreg_98 replaced by wreg_255

//ireg_92 replaced by ireg_239

//accumulate_99 replaced by accumulate_255

//umul_93 replaced by umul_239

//wreg_99 replaced by wreg_255

//ireg_93 replaced by ireg_239

//accumulate_100 replaced by accumulate_255

//umul_94 replaced by umul_239

//wreg_100 replaced by wreg_255

//ireg_94 replaced by ireg_239

//accumulate_101 replaced by accumulate_255

//umul_95 replaced by umul_239

//wreg_101 replaced by wreg_255

//ireg_95 replaced by ireg_239

//accumulate_102 replaced by accumulate_255

//umul_96 replaced by umul_239

//wreg_102 replaced by wreg_255

//ireg_96 replaced by ireg_239

//accumulate_103 replaced by accumulate_255

//umul_97 replaced by umul_239

//wreg_103 replaced by wreg_255

//ireg_97 replaced by ireg_239

//accumulate_104 replaced by accumulate_255

//umul_98 replaced by umul_239

//wreg_104 replaced by wreg_255

//ireg_98 replaced by ireg_239

//accumulate_105 replaced by accumulate_255

//umul_99 replaced by umul_239

//wreg_105 replaced by wreg_255

//ireg_99 replaced by ireg_239

//accumulate_106 replaced by accumulate_255

//umul_100 replaced by umul_239

//wreg_106 replaced by wreg_255

//ireg_100 replaced by ireg_239

//accumulate_107 replaced by accumulate_255

//umul_101 replaced by umul_239

//wreg_107 replaced by wreg_255

//ireg_101 replaced by ireg_239

//accumulate_108 replaced by accumulate_255

//umul_102 replaced by umul_239

//wreg_108 replaced by wreg_255

//ireg_102 replaced by ireg_239

//accumulate_109 replaced by accumulate_255

//umul_103 replaced by umul_239

//wreg_109 replaced by wreg_255

//ireg_103 replaced by ireg_239

//accumulate_110 replaced by accumulate_255

//umul_104 replaced by umul_239

//wreg_110 replaced by wreg_255

//ireg_104 replaced by ireg_239

//accumulate_111 replaced by accumulate_255

//umulBorder_6 replaced by umulBorder_15

//wreg_111 replaced by wreg_255

//uregBorder_6 replaced by uregBorder_15

//accumulate_112 replaced by accumulate_255

//umul_105 replaced by umul_239

//wreg_112 replaced by wreg_255

//ireg_105 replaced by ireg_239

//accumulate_113 replaced by accumulate_255

//umul_106 replaced by umul_239

//wreg_113 replaced by wreg_255

//ireg_106 replaced by ireg_239

//accumulate_114 replaced by accumulate_255

//umul_107 replaced by umul_239

//wreg_114 replaced by wreg_255

//ireg_107 replaced by ireg_239

//accumulate_115 replaced by accumulate_255

//umul_108 replaced by umul_239

//wreg_115 replaced by wreg_255

//ireg_108 replaced by ireg_239

//accumulate_116 replaced by accumulate_255

//umul_109 replaced by umul_239

//wreg_116 replaced by wreg_255

//ireg_109 replaced by ireg_239

//accumulate_117 replaced by accumulate_255

//umul_110 replaced by umul_239

//wreg_117 replaced by wreg_255

//ireg_110 replaced by ireg_239

//accumulate_118 replaced by accumulate_255

//umul_111 replaced by umul_239

//wreg_118 replaced by wreg_255

//ireg_111 replaced by ireg_239

//accumulate_119 replaced by accumulate_255

//umul_112 replaced by umul_239

//wreg_119 replaced by wreg_255

//ireg_112 replaced by ireg_239

//accumulate_120 replaced by accumulate_255

//umul_113 replaced by umul_239

//wreg_120 replaced by wreg_255

//ireg_113 replaced by ireg_239

//accumulate_121 replaced by accumulate_255

//umul_114 replaced by umul_239

//wreg_121 replaced by wreg_255

//ireg_114 replaced by ireg_239

//accumulate_122 replaced by accumulate_255

//umul_115 replaced by umul_239

//wreg_122 replaced by wreg_255

//ireg_115 replaced by ireg_239

//accumulate_123 replaced by accumulate_255

//umul_116 replaced by umul_239

//wreg_123 replaced by wreg_255

//ireg_116 replaced by ireg_239

//accumulate_124 replaced by accumulate_255

//umul_117 replaced by umul_239

//wreg_124 replaced by wreg_255

//ireg_117 replaced by ireg_239

//accumulate_125 replaced by accumulate_255

//umul_118 replaced by umul_239

//wreg_125 replaced by wreg_255

//ireg_118 replaced by ireg_239

//accumulate_126 replaced by accumulate_255

//umul_119 replaced by umul_239

//wreg_126 replaced by wreg_255

//ireg_119 replaced by ireg_239

//accumulate_127 replaced by accumulate_255

//umulBorder_7 replaced by umulBorder_15

//wreg_127 replaced by wreg_255

//uregBorder_7 replaced by uregBorder_15

//accumulate_128 replaced by accumulate_255

//umul_120 replaced by umul_239

//wreg_128 replaced by wreg_255

//ireg_120 replaced by ireg_239

//accumulate_129 replaced by accumulate_255

//umul_121 replaced by umul_239

//wreg_129 replaced by wreg_255

//ireg_121 replaced by ireg_239

//accumulate_130 replaced by accumulate_255

//umul_122 replaced by umul_239

//wreg_130 replaced by wreg_255

//ireg_122 replaced by ireg_239

//accumulate_131 replaced by accumulate_255

//umul_123 replaced by umul_239

//wreg_131 replaced by wreg_255

//ireg_123 replaced by ireg_239

//accumulate_132 replaced by accumulate_255

//umul_124 replaced by umul_239

//wreg_132 replaced by wreg_255

//ireg_124 replaced by ireg_239

//accumulate_133 replaced by accumulate_255

//umul_125 replaced by umul_239

//wreg_133 replaced by wreg_255

//ireg_125 replaced by ireg_239

//accumulate_134 replaced by accumulate_255

//umul_126 replaced by umul_239

//wreg_134 replaced by wreg_255

//ireg_126 replaced by ireg_239

//accumulate_135 replaced by accumulate_255

//umul_127 replaced by umul_239

//wreg_135 replaced by wreg_255

//ireg_127 replaced by ireg_239

//accumulate_136 replaced by accumulate_255

//umul_128 replaced by umul_239

//wreg_136 replaced by wreg_255

//ireg_128 replaced by ireg_239

//accumulate_137 replaced by accumulate_255

//umul_129 replaced by umul_239

//wreg_137 replaced by wreg_255

//ireg_129 replaced by ireg_239

//accumulate_138 replaced by accumulate_255

//umul_130 replaced by umul_239

//wreg_138 replaced by wreg_255

//ireg_130 replaced by ireg_239

//accumulate_139 replaced by accumulate_255

//umul_131 replaced by umul_239

//wreg_139 replaced by wreg_255

//ireg_131 replaced by ireg_239

//accumulate_140 replaced by accumulate_255

//umul_132 replaced by umul_239

//wreg_140 replaced by wreg_255

//ireg_132 replaced by ireg_239

//accumulate_141 replaced by accumulate_255

//umul_133 replaced by umul_239

//wreg_141 replaced by wreg_255

//ireg_133 replaced by ireg_239

//accumulate_142 replaced by accumulate_255

//umul_134 replaced by umul_239

//wreg_142 replaced by wreg_255

//ireg_134 replaced by ireg_239

//accumulate_143 replaced by accumulate_255

//umulBorder_8 replaced by umulBorder_15

//wreg_143 replaced by wreg_255

//uregBorder_8 replaced by uregBorder_15

//accumulate_144 replaced by accumulate_255

//umul_135 replaced by umul_239

//wreg_144 replaced by wreg_255

//ireg_135 replaced by ireg_239

//accumulate_145 replaced by accumulate_255

//umul_136 replaced by umul_239

//wreg_145 replaced by wreg_255

//ireg_136 replaced by ireg_239

//accumulate_146 replaced by accumulate_255

//umul_137 replaced by umul_239

//wreg_146 replaced by wreg_255

//ireg_137 replaced by ireg_239

//accumulate_147 replaced by accumulate_255

//umul_138 replaced by umul_239

//wreg_147 replaced by wreg_255

//ireg_138 replaced by ireg_239

//accumulate_148 replaced by accumulate_255

//umul_139 replaced by umul_239

//wreg_148 replaced by wreg_255

//ireg_139 replaced by ireg_239

//accumulate_149 replaced by accumulate_255

//umul_140 replaced by umul_239

//wreg_149 replaced by wreg_255

//ireg_140 replaced by ireg_239

//accumulate_150 replaced by accumulate_255

//umul_141 replaced by umul_239

//wreg_150 replaced by wreg_255

//ireg_141 replaced by ireg_239

//accumulate_151 replaced by accumulate_255

//umul_142 replaced by umul_239

//wreg_151 replaced by wreg_255

//ireg_142 replaced by ireg_239

//accumulate_152 replaced by accumulate_255

//umul_143 replaced by umul_239

//wreg_152 replaced by wreg_255

//ireg_143 replaced by ireg_239

//accumulate_153 replaced by accumulate_255

//umul_144 replaced by umul_239

//wreg_153 replaced by wreg_255

//ireg_144 replaced by ireg_239

//accumulate_154 replaced by accumulate_255

//umul_145 replaced by umul_239

//wreg_154 replaced by wreg_255

//ireg_145 replaced by ireg_239

//accumulate_155 replaced by accumulate_255

//umul_146 replaced by umul_239

//wreg_155 replaced by wreg_255

//ireg_146 replaced by ireg_239

//accumulate_156 replaced by accumulate_255

//umul_147 replaced by umul_239

//wreg_156 replaced by wreg_255

//ireg_147 replaced by ireg_239

//accumulate_157 replaced by accumulate_255

//umul_148 replaced by umul_239

//wreg_157 replaced by wreg_255

//ireg_148 replaced by ireg_239

//accumulate_158 replaced by accumulate_255

//umul_149 replaced by umul_239

//wreg_158 replaced by wreg_255

//ireg_149 replaced by ireg_239

//accumulate_159 replaced by accumulate_255

//umulBorder_9 replaced by umulBorder_15

//wreg_159 replaced by wreg_255

//uregBorder_9 replaced by uregBorder_15

//accumulate_160 replaced by accumulate_255

//umul_150 replaced by umul_239

//wreg_160 replaced by wreg_255

//ireg_150 replaced by ireg_239

//accumulate_161 replaced by accumulate_255

//umul_151 replaced by umul_239

//wreg_161 replaced by wreg_255

//ireg_151 replaced by ireg_239

//accumulate_162 replaced by accumulate_255

//umul_152 replaced by umul_239

//wreg_162 replaced by wreg_255

//ireg_152 replaced by ireg_239

//accumulate_163 replaced by accumulate_255

//umul_153 replaced by umul_239

//wreg_163 replaced by wreg_255

//ireg_153 replaced by ireg_239

//accumulate_164 replaced by accumulate_255

//umul_154 replaced by umul_239

//wreg_164 replaced by wreg_255

//ireg_154 replaced by ireg_239

//accumulate_165 replaced by accumulate_255

//umul_155 replaced by umul_239

//wreg_165 replaced by wreg_255

//ireg_155 replaced by ireg_239

//accumulate_166 replaced by accumulate_255

//umul_156 replaced by umul_239

//wreg_166 replaced by wreg_255

//ireg_156 replaced by ireg_239

//accumulate_167 replaced by accumulate_255

//umul_157 replaced by umul_239

//wreg_167 replaced by wreg_255

//ireg_157 replaced by ireg_239

//accumulate_168 replaced by accumulate_255

//umul_158 replaced by umul_239

//wreg_168 replaced by wreg_255

//ireg_158 replaced by ireg_239

//accumulate_169 replaced by accumulate_255

//umul_159 replaced by umul_239

//wreg_169 replaced by wreg_255

//ireg_159 replaced by ireg_239

//accumulate_170 replaced by accumulate_255

//umul_160 replaced by umul_239

//wreg_170 replaced by wreg_255

//ireg_160 replaced by ireg_239

//accumulate_171 replaced by accumulate_255

//umul_161 replaced by umul_239

//wreg_171 replaced by wreg_255

//ireg_161 replaced by ireg_239

//accumulate_172 replaced by accumulate_255

//umul_162 replaced by umul_239

//wreg_172 replaced by wreg_255

//ireg_162 replaced by ireg_239

//accumulate_173 replaced by accumulate_255

//umul_163 replaced by umul_239

//wreg_173 replaced by wreg_255

//ireg_163 replaced by ireg_239

//accumulate_174 replaced by accumulate_255

//umul_164 replaced by umul_239

//wreg_174 replaced by wreg_255

//ireg_164 replaced by ireg_239

//accumulate_175 replaced by accumulate_255

//umulBorder_10 replaced by umulBorder_15

//wreg_175 replaced by wreg_255

//uregBorder_10 replaced by uregBorder_15

//accumulate_176 replaced by accumulate_255

//umul_165 replaced by umul_239

//wreg_176 replaced by wreg_255

//ireg_165 replaced by ireg_239

//accumulate_177 replaced by accumulate_255

//umul_166 replaced by umul_239

//wreg_177 replaced by wreg_255

//ireg_166 replaced by ireg_239

//accumulate_178 replaced by accumulate_255

//umul_167 replaced by umul_239

//wreg_178 replaced by wreg_255

//ireg_167 replaced by ireg_239

//accumulate_179 replaced by accumulate_255

//umul_168 replaced by umul_239

//wreg_179 replaced by wreg_255

//ireg_168 replaced by ireg_239

//accumulate_180 replaced by accumulate_255

//umul_169 replaced by umul_239

//wreg_180 replaced by wreg_255

//ireg_169 replaced by ireg_239

//accumulate_181 replaced by accumulate_255

//umul_170 replaced by umul_239

//wreg_181 replaced by wreg_255

//ireg_170 replaced by ireg_239

//accumulate_182 replaced by accumulate_255

//umul_171 replaced by umul_239

//wreg_182 replaced by wreg_255

//ireg_171 replaced by ireg_239

//accumulate_183 replaced by accumulate_255

//umul_172 replaced by umul_239

//wreg_183 replaced by wreg_255

//ireg_172 replaced by ireg_239

//accumulate_184 replaced by accumulate_255

//umul_173 replaced by umul_239

//wreg_184 replaced by wreg_255

//ireg_173 replaced by ireg_239

//accumulate_185 replaced by accumulate_255

//umul_174 replaced by umul_239

//wreg_185 replaced by wreg_255

//ireg_174 replaced by ireg_239

//accumulate_186 replaced by accumulate_255

//umul_175 replaced by umul_239

//wreg_186 replaced by wreg_255

//ireg_175 replaced by ireg_239

//accumulate_187 replaced by accumulate_255

//umul_176 replaced by umul_239

//wreg_187 replaced by wreg_255

//ireg_176 replaced by ireg_239

//accumulate_188 replaced by accumulate_255

//umul_177 replaced by umul_239

//wreg_188 replaced by wreg_255

//ireg_177 replaced by ireg_239

//accumulate_189 replaced by accumulate_255

//umul_178 replaced by umul_239

//wreg_189 replaced by wreg_255

//ireg_178 replaced by ireg_239

//accumulate_190 replaced by accumulate_255

//umul_179 replaced by umul_239

//wreg_190 replaced by wreg_255

//ireg_179 replaced by ireg_239

//accumulate_191 replaced by accumulate_255

//umulBorder_11 replaced by umulBorder_15

//wreg_191 replaced by wreg_255

//uregBorder_11 replaced by uregBorder_15

//accumulate_192 replaced by accumulate_255

//umul_180 replaced by umul_239

//wreg_192 replaced by wreg_255

//ireg_180 replaced by ireg_239

//accumulate_193 replaced by accumulate_255

//umul_181 replaced by umul_239

//wreg_193 replaced by wreg_255

//ireg_181 replaced by ireg_239

//accumulate_194 replaced by accumulate_255

//umul_182 replaced by umul_239

//wreg_194 replaced by wreg_255

//ireg_182 replaced by ireg_239

//accumulate_195 replaced by accumulate_255

//umul_183 replaced by umul_239

//wreg_195 replaced by wreg_255

//ireg_183 replaced by ireg_239

//accumulate_196 replaced by accumulate_255

//umul_184 replaced by umul_239

//wreg_196 replaced by wreg_255

//ireg_184 replaced by ireg_239

//accumulate_197 replaced by accumulate_255

//umul_185 replaced by umul_239

//wreg_197 replaced by wreg_255

//ireg_185 replaced by ireg_239

//accumulate_198 replaced by accumulate_255

//umul_186 replaced by umul_239

//wreg_198 replaced by wreg_255

//ireg_186 replaced by ireg_239

//accumulate_199 replaced by accumulate_255

//umul_187 replaced by umul_239

//wreg_199 replaced by wreg_255

//ireg_187 replaced by ireg_239

//accumulate_200 replaced by accumulate_255

//umul_188 replaced by umul_239

//wreg_200 replaced by wreg_255

//ireg_188 replaced by ireg_239

//accumulate_201 replaced by accumulate_255

//umul_189 replaced by umul_239

//wreg_201 replaced by wreg_255

//ireg_189 replaced by ireg_239

//accumulate_202 replaced by accumulate_255

//umul_190 replaced by umul_239

//wreg_202 replaced by wreg_255

//ireg_190 replaced by ireg_239

//accumulate_203 replaced by accumulate_255

//umul_191 replaced by umul_239

//wreg_203 replaced by wreg_255

//ireg_191 replaced by ireg_239

//accumulate_204 replaced by accumulate_255

//umul_192 replaced by umul_239

//wreg_204 replaced by wreg_255

//ireg_192 replaced by ireg_239

//accumulate_205 replaced by accumulate_255

//umul_193 replaced by umul_239

//wreg_205 replaced by wreg_255

//ireg_193 replaced by ireg_239

//accumulate_206 replaced by accumulate_255

//umul_194 replaced by umul_239

//wreg_206 replaced by wreg_255

//ireg_194 replaced by ireg_239

//accumulate_207 replaced by accumulate_255

//umulBorder_12 replaced by umulBorder_15

//wreg_207 replaced by wreg_255

//uregBorder_12 replaced by uregBorder_15

//accumulate_208 replaced by accumulate_255

//umul_195 replaced by umul_239

//wreg_208 replaced by wreg_255

//ireg_195 replaced by ireg_239

//accumulate_209 replaced by accumulate_255

//umul_196 replaced by umul_239

//wreg_209 replaced by wreg_255

//ireg_196 replaced by ireg_239

//accumulate_210 replaced by accumulate_255

//umul_197 replaced by umul_239

//wreg_210 replaced by wreg_255

//ireg_197 replaced by ireg_239

//accumulate_211 replaced by accumulate_255

//umul_198 replaced by umul_239

//wreg_211 replaced by wreg_255

//ireg_198 replaced by ireg_239

//accumulate_212 replaced by accumulate_255

//umul_199 replaced by umul_239

//wreg_212 replaced by wreg_255

//ireg_199 replaced by ireg_239

//accumulate_213 replaced by accumulate_255

//umul_200 replaced by umul_239

//wreg_213 replaced by wreg_255

//ireg_200 replaced by ireg_239

//accumulate_214 replaced by accumulate_255

//umul_201 replaced by umul_239

//wreg_214 replaced by wreg_255

//ireg_201 replaced by ireg_239

//accumulate_215 replaced by accumulate_255

//umul_202 replaced by umul_239

//wreg_215 replaced by wreg_255

//ireg_202 replaced by ireg_239

//accumulate_216 replaced by accumulate_255

//umul_203 replaced by umul_239

//wreg_216 replaced by wreg_255

//ireg_203 replaced by ireg_239

//accumulate_217 replaced by accumulate_255

//umul_204 replaced by umul_239

//wreg_217 replaced by wreg_255

//ireg_204 replaced by ireg_239

//accumulate_218 replaced by accumulate_255

//umul_205 replaced by umul_239

//wreg_218 replaced by wreg_255

//ireg_205 replaced by ireg_239

//accumulate_219 replaced by accumulate_255

//umul_206 replaced by umul_239

//wreg_219 replaced by wreg_255

//ireg_206 replaced by ireg_239

//accumulate_220 replaced by accumulate_255

//umul_207 replaced by umul_239

//wreg_220 replaced by wreg_255

//ireg_207 replaced by ireg_239

//accumulate_221 replaced by accumulate_255

//umul_208 replaced by umul_239

//wreg_221 replaced by wreg_255

//ireg_208 replaced by ireg_239

//accumulate_222 replaced by accumulate_255

//umul_209 replaced by umul_239

//wreg_222 replaced by wreg_255

//ireg_209 replaced by ireg_239

//accumulate_223 replaced by accumulate_255

//umulBorder_13 replaced by umulBorder_15

//wreg_223 replaced by wreg_255

//uregBorder_13 replaced by uregBorder_15

//accumulate_224 replaced by accumulate_255

//umul_210 replaced by umul_239

//wreg_224 replaced by wreg_255

//ireg_210 replaced by ireg_239

//accumulate_225 replaced by accumulate_255

//umul_211 replaced by umul_239

//wreg_225 replaced by wreg_255

//ireg_211 replaced by ireg_239

//accumulate_226 replaced by accumulate_255

//umul_212 replaced by umul_239

//wreg_226 replaced by wreg_255

//ireg_212 replaced by ireg_239

//accumulate_227 replaced by accumulate_255

//umul_213 replaced by umul_239

//wreg_227 replaced by wreg_255

//ireg_213 replaced by ireg_239

//accumulate_228 replaced by accumulate_255

//umul_214 replaced by umul_239

//wreg_228 replaced by wreg_255

//ireg_214 replaced by ireg_239

//accumulate_229 replaced by accumulate_255

//umul_215 replaced by umul_239

//wreg_229 replaced by wreg_255

//ireg_215 replaced by ireg_239

//accumulate_230 replaced by accumulate_255

//umul_216 replaced by umul_239

//wreg_230 replaced by wreg_255

//ireg_216 replaced by ireg_239

//accumulate_231 replaced by accumulate_255

//umul_217 replaced by umul_239

//wreg_231 replaced by wreg_255

//ireg_217 replaced by ireg_239

//accumulate_232 replaced by accumulate_255

//umul_218 replaced by umul_239

//wreg_232 replaced by wreg_255

//ireg_218 replaced by ireg_239

//accumulate_233 replaced by accumulate_255

//umul_219 replaced by umul_239

//wreg_233 replaced by wreg_255

//ireg_219 replaced by ireg_239

//accumulate_234 replaced by accumulate_255

//umul_220 replaced by umul_239

//wreg_234 replaced by wreg_255

//ireg_220 replaced by ireg_239

//accumulate_235 replaced by accumulate_255

//umul_221 replaced by umul_239

//wreg_235 replaced by wreg_255

//ireg_221 replaced by ireg_239

//accumulate_236 replaced by accumulate_255

//umul_222 replaced by umul_239

//wreg_236 replaced by wreg_255

//ireg_222 replaced by ireg_239

//accumulate_237 replaced by accumulate_255

//umul_223 replaced by umul_239

//wreg_237 replaced by wreg_255

//ireg_223 replaced by ireg_239

//accumulate_238 replaced by accumulate_255

//umul_224 replaced by umul_239

//wreg_238 replaced by wreg_255

//ireg_224 replaced by ireg_239

//accumulate_239 replaced by accumulate_255

//umulBorder_14 replaced by umulBorder_15

//wreg_239 replaced by wreg_255

//uregBorder_14 replaced by uregBorder_15

//accumulate_240 replaced by accumulate_255

//umul_225 replaced by umul_239

//wreg_240 replaced by wreg_255

//ireg_225 replaced by ireg_239

//accumulate_241 replaced by accumulate_255

//umul_226 replaced by umul_239

//wreg_241 replaced by wreg_255

//ireg_226 replaced by ireg_239

//accumulate_242 replaced by accumulate_255

//umul_227 replaced by umul_239

//wreg_242 replaced by wreg_255

//ireg_227 replaced by ireg_239

//accumulate_243 replaced by accumulate_255

//umul_228 replaced by umul_239

//wreg_243 replaced by wreg_255

//ireg_228 replaced by ireg_239

//accumulate_244 replaced by accumulate_255

//umul_229 replaced by umul_239

//wreg_244 replaced by wreg_255

//ireg_229 replaced by ireg_239

//accumulate_245 replaced by accumulate_255

//umul_230 replaced by umul_239

//wreg_245 replaced by wreg_255

//ireg_230 replaced by ireg_239

//accumulate_246 replaced by accumulate_255

//umul_231 replaced by umul_239

//wreg_246 replaced by wreg_255

//ireg_231 replaced by ireg_239

//accumulate_247 replaced by accumulate_255

//umul_232 replaced by umul_239

//wreg_247 replaced by wreg_255

//ireg_232 replaced by ireg_239

//accumulate_248 replaced by accumulate_255

//umul_233 replaced by umul_239

//wreg_248 replaced by wreg_255

//ireg_233 replaced by ireg_239

//accumulate_249 replaced by accumulate_255

//umul_234 replaced by umul_239

//wreg_249 replaced by wreg_255

//ireg_234 replaced by ireg_239

//accumulate_250 replaced by accumulate_255

//umul_235 replaced by umul_239

//wreg_250 replaced by wreg_255

//ireg_235 replaced by ireg_239

//accumulate_251 replaced by accumulate_255

//umul_236 replaced by umul_239

//wreg_251 replaced by wreg_255

//ireg_236 replaced by ireg_239

//accumulate_252 replaced by accumulate_255

//umul_237 replaced by umul_239

//wreg_252 replaced by wreg_255

//ireg_237 replaced by ireg_239

//accumulate_253 replaced by accumulate_255

//umul_238 replaced by umul_239

//wreg_253 replaced by wreg_255

//ireg_238 replaced by ireg_239

//accumulate_254 replaced by accumulate_255

module umul_239 (
  input  wire          io_i_bit_i,
  input  wire [14:0]   io_i_data_w,
  input  wire [14:0]   io_i_randw,
  output wire [14:0]   io_o_randw,
  output wire          io_o_bit
);

  wire                bitW;

  assign bitW = (io_o_randw < io_i_data_w);
  assign io_o_bit = (io_i_bit_i && bitW);
  assign io_o_randw = io_i_randw;

endmodule

//wreg_254 replaced by wreg_255

module ireg_239 (
  input  wire          io_enable,
  input  wire          io_clear,
  input  wire          io_i_data_sign,
  input  wire          io_i_data_dff,
  output wire          io_o_data_sign,
  output wire          io_o_data_dff,
  input  wire          clk,
  input  wire          reset
);

  reg                 o_data_sign;
  reg                 o_data_dff;

  assign io_o_data_dff = o_data_dff;
  assign io_o_data_sign = o_data_sign;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      o_data_sign <= 1'b0;
      o_data_dff <= 1'b0;
    end else begin
      if(io_clear) begin
        o_data_dff <= 1'b0;
        o_data_sign <= 1'b0;
      end else begin
        if(io_enable) begin
          o_data_sign <= io_i_data_sign;
          o_data_dff <= io_i_data_dff;
        end
      end
    end
  end


endmodule

module accumulate_255 (
  input  wire          io_enable,
  input  wire          io_clear,
  input  wire          io_mac_done,
  input  wire          io_sign_activation,
  input  wire          io_sign_weight,
  input  wire [31:0]   io_sum_input,
  output wire [31:0]   io_sum_output,
  input  wire          io_prod_bit,
  input  wire          clk,
  input  wire          reset
);

  wire       [31:0]   _zz_prod;
  wire       [31:0]   _zz_sum_o;
  wire       [31:0]   _zz_sum_o_1;
  wire                neg;
  wire       [31:0]   prod;
  reg        [31:0]   sum_o;

  assign _zz_prod = (neg ? 32'hffffffff : 32'h00000001);
  assign _zz_sum_o = ($signed(io_sum_input) + $signed(sum_o));
  assign _zz_sum_o_1 = ($signed(sum_o) + $signed(prod));
  assign neg = (io_sign_weight ^ io_sign_activation);
  assign prod = (io_prod_bit ? _zz_prod : 32'h00000000);
  assign io_sum_output = sum_o;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      sum_o <= 32'h00000000;
    end else begin
      if(io_clear) begin
        sum_o <= 32'h00000000;
      end else begin
        if(io_enable) begin
          sum_o <= (io_mac_done ? _zz_sum_o : _zz_sum_o_1);
        end
      end
    end
  end


endmodule

module umulBorder_15 (
  input  wire          io_clear,
  input  wire          io_init,
  input  wire [14:0]   io_i_data_i,
  input  wire [14:0]   io_i_data_w,
  output wire [14:0]   io_randW,
  output wire          io_o_bit,
  output wire          io_i_bit_d,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   sobol_w_io_sobolSeq;
  reg        [14:0]   cnt;
  reg        [15:0]   randW_all;
  wire                bitI;
  wire                bitW;
  wire                o_bit;
  wire                when_umul_l41;

  sobol_15 sobol_w (
    .io_enable   (bitI                     ), //i
    .io_sobolSeq (sobol_w_io_sobolSeq[15:0]), //o
    .clk         (clk                      ), //i
    .reset       (reset                    )  //i
  );
  assign bitI = (! (cnt == 15'h0000));
  assign bitW = (io_randW < io_i_data_w);
  assign o_bit = (bitI && bitW);
  assign when_umul_l41 = (io_clear || (! bitI));
  assign io_randW = randW_all[15 : 1];
  assign io_o_bit = o_bit;
  assign io_i_bit_d = bitI;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      cnt <= 15'h0000;
      randW_all <= 16'h0000;
    end else begin
      if(io_init) begin
        cnt <= io_i_data_i;
      end else begin
        if(when_umul_l41) begin
          cnt <= 15'h0000;
        end else begin
          cnt <= (cnt - 15'h0001);
        end
      end
      randW_all <= sobol_w_io_sobolSeq;
    end
  end


endmodule

module wreg_255 (
  input  wire          io_enable,
  input  wire          io_clear,
  input  wire [14:0]   io_input_abs,
  input  wire          io_input_sign,
  output wire [14:0]   io_output_abs,
  output wire          io_output_sign,
  input  wire          clk,
  input  wire          reset
);

  reg        [14:0]   output_abs;
  reg                 output_sign;

  assign io_output_abs = output_abs;
  assign io_output_sign = output_sign;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      output_abs <= 15'h0000;
      output_sign <= 1'b0;
    end else begin
      if(io_clear) begin
        output_abs <= 15'h0000;
        output_sign <= 1'b0;
      end else begin
        if(io_enable) begin
          output_sign <= io_input_sign;
          output_abs <= io_input_abs;
        end
      end
    end
  end


endmodule

module uregBorder_15 (
  input  wire          io_enable,
  input  wire          io_clear,
  input  wire [15:0]   io_input,
  output wire          io_output_sign,
  output wire [14:0]   io_output_abs,
  input  wire          clk,
  input  wire          reset
);

  wire       [14:0]   _zz_io_output_abs;
  wire       [14:0]   _zz_io_output_abs_1;
  reg        [15:0]   output_data;
  wire       [15:0]   output_data_neg;

  assign _zz_io_output_abs = output_data_neg[14 : 0];
  assign _zz_io_output_abs_1 = output_data[14 : 0];
  assign output_data_neg = (- output_data);
  assign io_output_sign = output_data[15];
  assign io_output_abs = (io_output_sign ? _zz_io_output_abs : _zz_io_output_abs_1);
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      output_data <= 16'h0000;
    end else begin
      if(io_clear) begin
        output_data <= 16'h0000;
      end else begin
        if(io_enable) begin
          output_data <= io_input;
        end
      end
    end
  end


endmodule

//sobol replaced by sobol_15

//sobol_1 replaced by sobol_15

//sobol_2 replaced by sobol_15

//sobol_3 replaced by sobol_15

//sobol_4 replaced by sobol_15

//sobol_5 replaced by sobol_15

//sobol_6 replaced by sobol_15

//sobol_7 replaced by sobol_15

//sobol_8 replaced by sobol_15

//sobol_9 replaced by sobol_15

//sobol_10 replaced by sobol_15

//sobol_11 replaced by sobol_15

//sobol_12 replaced by sobol_15

//sobol_13 replaced by sobol_15

//sobol_14 replaced by sobol_15

module sobol_15 (
  input  wire          io_enable,
  output wire [15:0]   io_sobolSeq,
  input  wire          clk,
  input  wire          reset
);

  reg        [15:0]   _zz_sebolSeq;
  wire       [15:0]   dirvec_0;
  wire       [15:0]   dirvec_1;
  wire       [15:0]   dirvec_2;
  wire       [15:0]   dirvec_3;
  wire       [15:0]   dirvec_4;
  wire       [15:0]   dirvec_5;
  wire       [15:0]   dirvec_6;
  wire       [15:0]   dirvec_7;
  wire       [15:0]   dirvec_8;
  wire       [15:0]   dirvec_9;
  wire       [15:0]   dirvec_10;
  wire       [15:0]   dirvec_11;
  wire       [15:0]   dirvec_12;
  wire       [15:0]   dirvec_13;
  wire       [15:0]   dirvec_14;
  wire       [15:0]   dirvec_15;
  reg        [3:0]    vecIdx;
  reg        [15:0]   cnt;
  reg        [15:0]   inacc;
  reg        [15:0]   outoh;
  reg        [15:0]   sebolSeq;

  always @(*) begin
    case(vecIdx)
      4'b0000 : _zz_sebolSeq = dirvec_0;
      4'b0001 : _zz_sebolSeq = dirvec_1;
      4'b0010 : _zz_sebolSeq = dirvec_2;
      4'b0011 : _zz_sebolSeq = dirvec_3;
      4'b0100 : _zz_sebolSeq = dirvec_4;
      4'b0101 : _zz_sebolSeq = dirvec_5;
      4'b0110 : _zz_sebolSeq = dirvec_6;
      4'b0111 : _zz_sebolSeq = dirvec_7;
      4'b1000 : _zz_sebolSeq = dirvec_8;
      4'b1001 : _zz_sebolSeq = dirvec_9;
      4'b1010 : _zz_sebolSeq = dirvec_10;
      4'b1011 : _zz_sebolSeq = dirvec_11;
      4'b1100 : _zz_sebolSeq = dirvec_12;
      4'b1101 : _zz_sebolSeq = dirvec_13;
      4'b1110 : _zz_sebolSeq = dirvec_14;
      default : _zz_sebolSeq = dirvec_15;
    endcase
  end

  always @(*) begin
    inacc[0] = (! cnt[0]);
    inacc[1] = (inacc[0] || (! cnt[1]));
    inacc[2] = (inacc[1] || (! cnt[2]));
    inacc[3] = (inacc[2] || (! cnt[3]));
    inacc[4] = (inacc[3] || (! cnt[4]));
    inacc[5] = (inacc[4] || (! cnt[5]));
    inacc[6] = (inacc[5] || (! cnt[6]));
    inacc[7] = (inacc[6] || (! cnt[7]));
    inacc[8] = (inacc[7] || (! cnt[8]));
    inacc[9] = (inacc[8] || (! cnt[9]));
    inacc[10] = (inacc[9] || (! cnt[10]));
    inacc[11] = (inacc[10] || (! cnt[11]));
    inacc[12] = (inacc[11] || (! cnt[12]));
    inacc[13] = (inacc[12] || (! cnt[13]));
    inacc[14] = (inacc[13] || (! cnt[14]));
    inacc[15] = (inacc[14] || (! cnt[15]));
  end

  always @(*) begin
    outoh[0] = (! cnt[0]);
    outoh[1] = (inacc[0] ^ inacc[1]);
    outoh[2] = (inacc[1] ^ inacc[2]);
    outoh[3] = (inacc[2] ^ inacc[3]);
    outoh[4] = (inacc[3] ^ inacc[4]);
    outoh[5] = (inacc[4] ^ inacc[5]);
    outoh[6] = (inacc[5] ^ inacc[6]);
    outoh[7] = (inacc[6] ^ inacc[7]);
    outoh[8] = (inacc[7] ^ inacc[8]);
    outoh[9] = (inacc[8] ^ inacc[9]);
    outoh[10] = (inacc[9] ^ inacc[10]);
    outoh[11] = (inacc[10] ^ inacc[11]);
    outoh[12] = (inacc[11] ^ inacc[12]);
    outoh[13] = (inacc[12] ^ inacc[13]);
    outoh[14] = (inacc[13] ^ inacc[14]);
    outoh[15] = (inacc[14] ^ inacc[15]);
  end

  assign dirvec_0 = 16'h8000;
  assign dirvec_1 = 16'h4000;
  assign dirvec_2 = 16'h2000;
  assign dirvec_3 = 16'h1000;
  assign dirvec_4 = 16'h0800;
  assign dirvec_5 = 16'h0400;
  assign dirvec_6 = 16'h0200;
  assign dirvec_7 = 16'h0100;
  assign dirvec_8 = 16'h0080;
  assign dirvec_9 = 16'h0040;
  assign dirvec_10 = 16'h0020;
  assign dirvec_11 = 16'h0010;
  assign dirvec_12 = 16'h0008;
  assign dirvec_13 = 16'h0004;
  assign dirvec_14 = 16'h0002;
  assign dirvec_15 = 16'h0001;
  always @(*) begin
    case(outoh)
      16'h0001 : begin
        vecIdx = 4'b0000;
      end
      16'h0002 : begin
        vecIdx = 4'b0001;
      end
      16'h0004 : begin
        vecIdx = 4'b0010;
      end
      16'h0008 : begin
        vecIdx = 4'b0011;
      end
      16'h0010 : begin
        vecIdx = 4'b0100;
      end
      16'h0020 : begin
        vecIdx = 4'b0101;
      end
      16'h0040 : begin
        vecIdx = 4'b0110;
      end
      16'h0080 : begin
        vecIdx = 4'b0111;
      end
      16'h0100 : begin
        vecIdx = 4'b1000;
      end
      16'h0200 : begin
        vecIdx = 4'b1001;
      end
      16'h0400 : begin
        vecIdx = 4'b1010;
      end
      16'h0800 : begin
        vecIdx = 4'b1011;
      end
      16'h1000 : begin
        vecIdx = 4'b1100;
      end
      16'h2000 : begin
        vecIdx = 4'b1101;
      end
      16'h4000 : begin
        vecIdx = 4'b1110;
      end
      16'h8000 : begin
        vecIdx = 4'b1111;
      end
      default : begin
        vecIdx = 4'b0000;
      end
    endcase
  end

  assign io_sobolSeq = sebolSeq;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      cnt <= 16'h0000;
      sebolSeq <= 16'h0000;
    end else begin
      if(io_enable) begin
        cnt <= (cnt + 16'h0001);
      end
      if(io_enable) begin
        sebolSeq <= (sebolSeq ^ _zz_sebolSeq);
      end
    end
  end


endmodule
