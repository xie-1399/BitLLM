// Generator : SpinalHDL v1.9.4    git head : 270018552577f3bb8e5339ee2583c9c22d324215
// Component : SystolicArray
// Git hash  : 95d4b99c2c5c0c9e41b84111df30141758565e63

`timescale 1ns/1ps

module SystolicArray (
  input  wire          io_load,
  input  wire [7:0]    io_activation_0,
  input  wire [7:0]    io_activation_1,
  input  wire [7:0]    io_activation_2,
  input  wire [7:0]    io_activation_3,
  input  wire [7:0]    io_activation_4,
  input  wire [7:0]    io_activation_5,
  input  wire [7:0]    io_activation_6,
  input  wire [7:0]    io_activation_7,
  input  wire [7:0]    io_activation_8,
  input  wire [7:0]    io_activation_9,
  input  wire [7:0]    io_activation_10,
  input  wire [7:0]    io_activation_11,
  input  wire [7:0]    io_activation_12,
  input  wire [7:0]    io_activation_13,
  input  wire [7:0]    io_activation_14,
  input  wire [7:0]    io_activation_15,
  input  wire [7:0]    io_activation_16,
  input  wire [7:0]    io_activation_17,
  input  wire [7:0]    io_activation_18,
  input  wire [7:0]    io_activation_19,
  input  wire [7:0]    io_activation_20,
  input  wire [7:0]    io_activation_21,
  input  wire [7:0]    io_activation_22,
  input  wire [7:0]    io_activation_23,
  input  wire [7:0]    io_activation_24,
  input  wire [7:0]    io_activation_25,
  input  wire [7:0]    io_activation_26,
  input  wire [7:0]    io_activation_27,
  input  wire [7:0]    io_activation_28,
  input  wire [7:0]    io_activation_29,
  input  wire [7:0]    io_activation_30,
  input  wire [7:0]    io_activation_31,
  input  wire [7:0]    io_weight_0,
  input  wire [7:0]    io_weight_1,
  input  wire [7:0]    io_weight_2,
  input  wire [7:0]    io_weight_3,
  input  wire [7:0]    io_weight_4,
  input  wire [7:0]    io_weight_5,
  input  wire [7:0]    io_weight_6,
  input  wire [7:0]    io_weight_7,
  input  wire [7:0]    io_weight_8,
  input  wire [7:0]    io_weight_9,
  input  wire [7:0]    io_weight_10,
  input  wire [7:0]    io_weight_11,
  input  wire [7:0]    io_weight_12,
  input  wire [7:0]    io_weight_13,
  input  wire [7:0]    io_weight_14,
  input  wire [7:0]    io_weight_15,
  input  wire [7:0]    io_weight_16,
  input  wire [7:0]    io_weight_17,
  input  wire [7:0]    io_weight_18,
  input  wire [7:0]    io_weight_19,
  input  wire [7:0]    io_weight_20,
  input  wire [7:0]    io_weight_21,
  input  wire [7:0]    io_weight_22,
  input  wire [7:0]    io_weight_23,
  input  wire [7:0]    io_weight_24,
  input  wire [7:0]    io_weight_25,
  input  wire [7:0]    io_weight_26,
  input  wire [7:0]    io_weight_27,
  input  wire [7:0]    io_weight_28,
  input  wire [7:0]    io_weight_29,
  input  wire [7:0]    io_weight_30,
  input  wire [7:0]    io_weight_31,
  output wire [7:0]    io_output_0,
  output wire [7:0]    io_output_1,
  output wire [7:0]    io_output_2,
  output wire [7:0]    io_output_3,
  output wire [7:0]    io_output_4,
  output wire [7:0]    io_output_5,
  output wire [7:0]    io_output_6,
  output wire [7:0]    io_output_7,
  output wire [7:0]    io_output_8,
  output wire [7:0]    io_output_9,
  output wire [7:0]    io_output_10,
  output wire [7:0]    io_output_11,
  output wire [7:0]    io_output_12,
  output wire [7:0]    io_output_13,
  output wire [7:0]    io_output_14,
  output wire [7:0]    io_output_15,
  output wire [7:0]    io_output_16,
  output wire [7:0]    io_output_17,
  output wire [7:0]    io_output_18,
  output wire [7:0]    io_output_19,
  output wire [7:0]    io_output_20,
  output wire [7:0]    io_output_21,
  output wire [7:0]    io_output_22,
  output wire [7:0]    io_output_23,
  output wire [7:0]    io_output_24,
  output wire [7:0]    io_output_25,
  output wire [7:0]    io_output_26,
  output wire [7:0]    io_output_27,
  output wire [7:0]    io_output_28,
  output wire [7:0]    io_output_29,
  output wire [7:0]    io_output_30,
  output wire [7:0]    io_output_31,
  input  wire          clk,
  input  wire          reset
);

  wire       [7:0]    mac_0_0_io_passthrough;
  wire       [7:0]    mac_0_0_io_macOut;
  wire       [7:0]    mac_0_1_io_passthrough;
  wire       [7:0]    mac_0_1_io_macOut;
  wire       [7:0]    mac_0_2_io_passthrough;
  wire       [7:0]    mac_0_2_io_macOut;
  wire       [7:0]    mac_0_3_io_passthrough;
  wire       [7:0]    mac_0_3_io_macOut;
  wire       [7:0]    mac_0_4_io_passthrough;
  wire       [7:0]    mac_0_4_io_macOut;
  wire       [7:0]    mac_0_5_io_passthrough;
  wire       [7:0]    mac_0_5_io_macOut;
  wire       [7:0]    mac_0_6_io_passthrough;
  wire       [7:0]    mac_0_6_io_macOut;
  wire       [7:0]    mac_0_7_io_passthrough;
  wire       [7:0]    mac_0_7_io_macOut;
  wire       [7:0]    mac_0_8_io_passthrough;
  wire       [7:0]    mac_0_8_io_macOut;
  wire       [7:0]    mac_0_9_io_passthrough;
  wire       [7:0]    mac_0_9_io_macOut;
  wire       [7:0]    mac_0_10_io_passthrough;
  wire       [7:0]    mac_0_10_io_macOut;
  wire       [7:0]    mac_0_11_io_passthrough;
  wire       [7:0]    mac_0_11_io_macOut;
  wire       [7:0]    mac_0_12_io_passthrough;
  wire       [7:0]    mac_0_12_io_macOut;
  wire       [7:0]    mac_0_13_io_passthrough;
  wire       [7:0]    mac_0_13_io_macOut;
  wire       [7:0]    mac_0_14_io_passthrough;
  wire       [7:0]    mac_0_14_io_macOut;
  wire       [7:0]    mac_0_15_io_passthrough;
  wire       [7:0]    mac_0_15_io_macOut;
  wire       [7:0]    mac_0_16_io_passthrough;
  wire       [7:0]    mac_0_16_io_macOut;
  wire       [7:0]    mac_0_17_io_passthrough;
  wire       [7:0]    mac_0_17_io_macOut;
  wire       [7:0]    mac_0_18_io_passthrough;
  wire       [7:0]    mac_0_18_io_macOut;
  wire       [7:0]    mac_0_19_io_passthrough;
  wire       [7:0]    mac_0_19_io_macOut;
  wire       [7:0]    mac_0_20_io_passthrough;
  wire       [7:0]    mac_0_20_io_macOut;
  wire       [7:0]    mac_0_21_io_passthrough;
  wire       [7:0]    mac_0_21_io_macOut;
  wire       [7:0]    mac_0_22_io_passthrough;
  wire       [7:0]    mac_0_22_io_macOut;
  wire       [7:0]    mac_0_23_io_passthrough;
  wire       [7:0]    mac_0_23_io_macOut;
  wire       [7:0]    mac_0_24_io_passthrough;
  wire       [7:0]    mac_0_24_io_macOut;
  wire       [7:0]    mac_0_25_io_passthrough;
  wire       [7:0]    mac_0_25_io_macOut;
  wire       [7:0]    mac_0_26_io_passthrough;
  wire       [7:0]    mac_0_26_io_macOut;
  wire       [7:0]    mac_0_27_io_passthrough;
  wire       [7:0]    mac_0_27_io_macOut;
  wire       [7:0]    mac_0_28_io_passthrough;
  wire       [7:0]    mac_0_28_io_macOut;
  wire       [7:0]    mac_0_29_io_passthrough;
  wire       [7:0]    mac_0_29_io_macOut;
  wire       [7:0]    mac_0_30_io_passthrough;
  wire       [7:0]    mac_0_30_io_macOut;
  wire       [7:0]    mac_0_31_io_passthrough;
  wire       [7:0]    mac_0_31_io_macOut;
  wire       [7:0]    mac_1_0_io_passthrough;
  wire       [7:0]    mac_1_0_io_macOut;
  wire       [7:0]    mac_1_1_io_passthrough;
  wire       [7:0]    mac_1_1_io_macOut;
  wire       [7:0]    mac_1_2_io_passthrough;
  wire       [7:0]    mac_1_2_io_macOut;
  wire       [7:0]    mac_1_3_io_passthrough;
  wire       [7:0]    mac_1_3_io_macOut;
  wire       [7:0]    mac_1_4_io_passthrough;
  wire       [7:0]    mac_1_4_io_macOut;
  wire       [7:0]    mac_1_5_io_passthrough;
  wire       [7:0]    mac_1_5_io_macOut;
  wire       [7:0]    mac_1_6_io_passthrough;
  wire       [7:0]    mac_1_6_io_macOut;
  wire       [7:0]    mac_1_7_io_passthrough;
  wire       [7:0]    mac_1_7_io_macOut;
  wire       [7:0]    mac_1_8_io_passthrough;
  wire       [7:0]    mac_1_8_io_macOut;
  wire       [7:0]    mac_1_9_io_passthrough;
  wire       [7:0]    mac_1_9_io_macOut;
  wire       [7:0]    mac_1_10_io_passthrough;
  wire       [7:0]    mac_1_10_io_macOut;
  wire       [7:0]    mac_1_11_io_passthrough;
  wire       [7:0]    mac_1_11_io_macOut;
  wire       [7:0]    mac_1_12_io_passthrough;
  wire       [7:0]    mac_1_12_io_macOut;
  wire       [7:0]    mac_1_13_io_passthrough;
  wire       [7:0]    mac_1_13_io_macOut;
  wire       [7:0]    mac_1_14_io_passthrough;
  wire       [7:0]    mac_1_14_io_macOut;
  wire       [7:0]    mac_1_15_io_passthrough;
  wire       [7:0]    mac_1_15_io_macOut;
  wire       [7:0]    mac_1_16_io_passthrough;
  wire       [7:0]    mac_1_16_io_macOut;
  wire       [7:0]    mac_1_17_io_passthrough;
  wire       [7:0]    mac_1_17_io_macOut;
  wire       [7:0]    mac_1_18_io_passthrough;
  wire       [7:0]    mac_1_18_io_macOut;
  wire       [7:0]    mac_1_19_io_passthrough;
  wire       [7:0]    mac_1_19_io_macOut;
  wire       [7:0]    mac_1_20_io_passthrough;
  wire       [7:0]    mac_1_20_io_macOut;
  wire       [7:0]    mac_1_21_io_passthrough;
  wire       [7:0]    mac_1_21_io_macOut;
  wire       [7:0]    mac_1_22_io_passthrough;
  wire       [7:0]    mac_1_22_io_macOut;
  wire       [7:0]    mac_1_23_io_passthrough;
  wire       [7:0]    mac_1_23_io_macOut;
  wire       [7:0]    mac_1_24_io_passthrough;
  wire       [7:0]    mac_1_24_io_macOut;
  wire       [7:0]    mac_1_25_io_passthrough;
  wire       [7:0]    mac_1_25_io_macOut;
  wire       [7:0]    mac_1_26_io_passthrough;
  wire       [7:0]    mac_1_26_io_macOut;
  wire       [7:0]    mac_1_27_io_passthrough;
  wire       [7:0]    mac_1_27_io_macOut;
  wire       [7:0]    mac_1_28_io_passthrough;
  wire       [7:0]    mac_1_28_io_macOut;
  wire       [7:0]    mac_1_29_io_passthrough;
  wire       [7:0]    mac_1_29_io_macOut;
  wire       [7:0]    mac_1_30_io_passthrough;
  wire       [7:0]    mac_1_30_io_macOut;
  wire       [7:0]    mac_1_31_io_passthrough;
  wire       [7:0]    mac_1_31_io_macOut;
  wire       [7:0]    mac_2_0_io_passthrough;
  wire       [7:0]    mac_2_0_io_macOut;
  wire       [7:0]    mac_2_1_io_passthrough;
  wire       [7:0]    mac_2_1_io_macOut;
  wire       [7:0]    mac_2_2_io_passthrough;
  wire       [7:0]    mac_2_2_io_macOut;
  wire       [7:0]    mac_2_3_io_passthrough;
  wire       [7:0]    mac_2_3_io_macOut;
  wire       [7:0]    mac_2_4_io_passthrough;
  wire       [7:0]    mac_2_4_io_macOut;
  wire       [7:0]    mac_2_5_io_passthrough;
  wire       [7:0]    mac_2_5_io_macOut;
  wire       [7:0]    mac_2_6_io_passthrough;
  wire       [7:0]    mac_2_6_io_macOut;
  wire       [7:0]    mac_2_7_io_passthrough;
  wire       [7:0]    mac_2_7_io_macOut;
  wire       [7:0]    mac_2_8_io_passthrough;
  wire       [7:0]    mac_2_8_io_macOut;
  wire       [7:0]    mac_2_9_io_passthrough;
  wire       [7:0]    mac_2_9_io_macOut;
  wire       [7:0]    mac_2_10_io_passthrough;
  wire       [7:0]    mac_2_10_io_macOut;
  wire       [7:0]    mac_2_11_io_passthrough;
  wire       [7:0]    mac_2_11_io_macOut;
  wire       [7:0]    mac_2_12_io_passthrough;
  wire       [7:0]    mac_2_12_io_macOut;
  wire       [7:0]    mac_2_13_io_passthrough;
  wire       [7:0]    mac_2_13_io_macOut;
  wire       [7:0]    mac_2_14_io_passthrough;
  wire       [7:0]    mac_2_14_io_macOut;
  wire       [7:0]    mac_2_15_io_passthrough;
  wire       [7:0]    mac_2_15_io_macOut;
  wire       [7:0]    mac_2_16_io_passthrough;
  wire       [7:0]    mac_2_16_io_macOut;
  wire       [7:0]    mac_2_17_io_passthrough;
  wire       [7:0]    mac_2_17_io_macOut;
  wire       [7:0]    mac_2_18_io_passthrough;
  wire       [7:0]    mac_2_18_io_macOut;
  wire       [7:0]    mac_2_19_io_passthrough;
  wire       [7:0]    mac_2_19_io_macOut;
  wire       [7:0]    mac_2_20_io_passthrough;
  wire       [7:0]    mac_2_20_io_macOut;
  wire       [7:0]    mac_2_21_io_passthrough;
  wire       [7:0]    mac_2_21_io_macOut;
  wire       [7:0]    mac_2_22_io_passthrough;
  wire       [7:0]    mac_2_22_io_macOut;
  wire       [7:0]    mac_2_23_io_passthrough;
  wire       [7:0]    mac_2_23_io_macOut;
  wire       [7:0]    mac_2_24_io_passthrough;
  wire       [7:0]    mac_2_24_io_macOut;
  wire       [7:0]    mac_2_25_io_passthrough;
  wire       [7:0]    mac_2_25_io_macOut;
  wire       [7:0]    mac_2_26_io_passthrough;
  wire       [7:0]    mac_2_26_io_macOut;
  wire       [7:0]    mac_2_27_io_passthrough;
  wire       [7:0]    mac_2_27_io_macOut;
  wire       [7:0]    mac_2_28_io_passthrough;
  wire       [7:0]    mac_2_28_io_macOut;
  wire       [7:0]    mac_2_29_io_passthrough;
  wire       [7:0]    mac_2_29_io_macOut;
  wire       [7:0]    mac_2_30_io_passthrough;
  wire       [7:0]    mac_2_30_io_macOut;
  wire       [7:0]    mac_2_31_io_passthrough;
  wire       [7:0]    mac_2_31_io_macOut;
  wire       [7:0]    mac_3_0_io_passthrough;
  wire       [7:0]    mac_3_0_io_macOut;
  wire       [7:0]    mac_3_1_io_passthrough;
  wire       [7:0]    mac_3_1_io_macOut;
  wire       [7:0]    mac_3_2_io_passthrough;
  wire       [7:0]    mac_3_2_io_macOut;
  wire       [7:0]    mac_3_3_io_passthrough;
  wire       [7:0]    mac_3_3_io_macOut;
  wire       [7:0]    mac_3_4_io_passthrough;
  wire       [7:0]    mac_3_4_io_macOut;
  wire       [7:0]    mac_3_5_io_passthrough;
  wire       [7:0]    mac_3_5_io_macOut;
  wire       [7:0]    mac_3_6_io_passthrough;
  wire       [7:0]    mac_3_6_io_macOut;
  wire       [7:0]    mac_3_7_io_passthrough;
  wire       [7:0]    mac_3_7_io_macOut;
  wire       [7:0]    mac_3_8_io_passthrough;
  wire       [7:0]    mac_3_8_io_macOut;
  wire       [7:0]    mac_3_9_io_passthrough;
  wire       [7:0]    mac_3_9_io_macOut;
  wire       [7:0]    mac_3_10_io_passthrough;
  wire       [7:0]    mac_3_10_io_macOut;
  wire       [7:0]    mac_3_11_io_passthrough;
  wire       [7:0]    mac_3_11_io_macOut;
  wire       [7:0]    mac_3_12_io_passthrough;
  wire       [7:0]    mac_3_12_io_macOut;
  wire       [7:0]    mac_3_13_io_passthrough;
  wire       [7:0]    mac_3_13_io_macOut;
  wire       [7:0]    mac_3_14_io_passthrough;
  wire       [7:0]    mac_3_14_io_macOut;
  wire       [7:0]    mac_3_15_io_passthrough;
  wire       [7:0]    mac_3_15_io_macOut;
  wire       [7:0]    mac_3_16_io_passthrough;
  wire       [7:0]    mac_3_16_io_macOut;
  wire       [7:0]    mac_3_17_io_passthrough;
  wire       [7:0]    mac_3_17_io_macOut;
  wire       [7:0]    mac_3_18_io_passthrough;
  wire       [7:0]    mac_3_18_io_macOut;
  wire       [7:0]    mac_3_19_io_passthrough;
  wire       [7:0]    mac_3_19_io_macOut;
  wire       [7:0]    mac_3_20_io_passthrough;
  wire       [7:0]    mac_3_20_io_macOut;
  wire       [7:0]    mac_3_21_io_passthrough;
  wire       [7:0]    mac_3_21_io_macOut;
  wire       [7:0]    mac_3_22_io_passthrough;
  wire       [7:0]    mac_3_22_io_macOut;
  wire       [7:0]    mac_3_23_io_passthrough;
  wire       [7:0]    mac_3_23_io_macOut;
  wire       [7:0]    mac_3_24_io_passthrough;
  wire       [7:0]    mac_3_24_io_macOut;
  wire       [7:0]    mac_3_25_io_passthrough;
  wire       [7:0]    mac_3_25_io_macOut;
  wire       [7:0]    mac_3_26_io_passthrough;
  wire       [7:0]    mac_3_26_io_macOut;
  wire       [7:0]    mac_3_27_io_passthrough;
  wire       [7:0]    mac_3_27_io_macOut;
  wire       [7:0]    mac_3_28_io_passthrough;
  wire       [7:0]    mac_3_28_io_macOut;
  wire       [7:0]    mac_3_29_io_passthrough;
  wire       [7:0]    mac_3_29_io_macOut;
  wire       [7:0]    mac_3_30_io_passthrough;
  wire       [7:0]    mac_3_30_io_macOut;
  wire       [7:0]    mac_3_31_io_passthrough;
  wire       [7:0]    mac_3_31_io_macOut;
  wire       [7:0]    mac_4_0_io_passthrough;
  wire       [7:0]    mac_4_0_io_macOut;
  wire       [7:0]    mac_4_1_io_passthrough;
  wire       [7:0]    mac_4_1_io_macOut;
  wire       [7:0]    mac_4_2_io_passthrough;
  wire       [7:0]    mac_4_2_io_macOut;
  wire       [7:0]    mac_4_3_io_passthrough;
  wire       [7:0]    mac_4_3_io_macOut;
  wire       [7:0]    mac_4_4_io_passthrough;
  wire       [7:0]    mac_4_4_io_macOut;
  wire       [7:0]    mac_4_5_io_passthrough;
  wire       [7:0]    mac_4_5_io_macOut;
  wire       [7:0]    mac_4_6_io_passthrough;
  wire       [7:0]    mac_4_6_io_macOut;
  wire       [7:0]    mac_4_7_io_passthrough;
  wire       [7:0]    mac_4_7_io_macOut;
  wire       [7:0]    mac_4_8_io_passthrough;
  wire       [7:0]    mac_4_8_io_macOut;
  wire       [7:0]    mac_4_9_io_passthrough;
  wire       [7:0]    mac_4_9_io_macOut;
  wire       [7:0]    mac_4_10_io_passthrough;
  wire       [7:0]    mac_4_10_io_macOut;
  wire       [7:0]    mac_4_11_io_passthrough;
  wire       [7:0]    mac_4_11_io_macOut;
  wire       [7:0]    mac_4_12_io_passthrough;
  wire       [7:0]    mac_4_12_io_macOut;
  wire       [7:0]    mac_4_13_io_passthrough;
  wire       [7:0]    mac_4_13_io_macOut;
  wire       [7:0]    mac_4_14_io_passthrough;
  wire       [7:0]    mac_4_14_io_macOut;
  wire       [7:0]    mac_4_15_io_passthrough;
  wire       [7:0]    mac_4_15_io_macOut;
  wire       [7:0]    mac_4_16_io_passthrough;
  wire       [7:0]    mac_4_16_io_macOut;
  wire       [7:0]    mac_4_17_io_passthrough;
  wire       [7:0]    mac_4_17_io_macOut;
  wire       [7:0]    mac_4_18_io_passthrough;
  wire       [7:0]    mac_4_18_io_macOut;
  wire       [7:0]    mac_4_19_io_passthrough;
  wire       [7:0]    mac_4_19_io_macOut;
  wire       [7:0]    mac_4_20_io_passthrough;
  wire       [7:0]    mac_4_20_io_macOut;
  wire       [7:0]    mac_4_21_io_passthrough;
  wire       [7:0]    mac_4_21_io_macOut;
  wire       [7:0]    mac_4_22_io_passthrough;
  wire       [7:0]    mac_4_22_io_macOut;
  wire       [7:0]    mac_4_23_io_passthrough;
  wire       [7:0]    mac_4_23_io_macOut;
  wire       [7:0]    mac_4_24_io_passthrough;
  wire       [7:0]    mac_4_24_io_macOut;
  wire       [7:0]    mac_4_25_io_passthrough;
  wire       [7:0]    mac_4_25_io_macOut;
  wire       [7:0]    mac_4_26_io_passthrough;
  wire       [7:0]    mac_4_26_io_macOut;
  wire       [7:0]    mac_4_27_io_passthrough;
  wire       [7:0]    mac_4_27_io_macOut;
  wire       [7:0]    mac_4_28_io_passthrough;
  wire       [7:0]    mac_4_28_io_macOut;
  wire       [7:0]    mac_4_29_io_passthrough;
  wire       [7:0]    mac_4_29_io_macOut;
  wire       [7:0]    mac_4_30_io_passthrough;
  wire       [7:0]    mac_4_30_io_macOut;
  wire       [7:0]    mac_4_31_io_passthrough;
  wire       [7:0]    mac_4_31_io_macOut;
  wire       [7:0]    mac_5_0_io_passthrough;
  wire       [7:0]    mac_5_0_io_macOut;
  wire       [7:0]    mac_5_1_io_passthrough;
  wire       [7:0]    mac_5_1_io_macOut;
  wire       [7:0]    mac_5_2_io_passthrough;
  wire       [7:0]    mac_5_2_io_macOut;
  wire       [7:0]    mac_5_3_io_passthrough;
  wire       [7:0]    mac_5_3_io_macOut;
  wire       [7:0]    mac_5_4_io_passthrough;
  wire       [7:0]    mac_5_4_io_macOut;
  wire       [7:0]    mac_5_5_io_passthrough;
  wire       [7:0]    mac_5_5_io_macOut;
  wire       [7:0]    mac_5_6_io_passthrough;
  wire       [7:0]    mac_5_6_io_macOut;
  wire       [7:0]    mac_5_7_io_passthrough;
  wire       [7:0]    mac_5_7_io_macOut;
  wire       [7:0]    mac_5_8_io_passthrough;
  wire       [7:0]    mac_5_8_io_macOut;
  wire       [7:0]    mac_5_9_io_passthrough;
  wire       [7:0]    mac_5_9_io_macOut;
  wire       [7:0]    mac_5_10_io_passthrough;
  wire       [7:0]    mac_5_10_io_macOut;
  wire       [7:0]    mac_5_11_io_passthrough;
  wire       [7:0]    mac_5_11_io_macOut;
  wire       [7:0]    mac_5_12_io_passthrough;
  wire       [7:0]    mac_5_12_io_macOut;
  wire       [7:0]    mac_5_13_io_passthrough;
  wire       [7:0]    mac_5_13_io_macOut;
  wire       [7:0]    mac_5_14_io_passthrough;
  wire       [7:0]    mac_5_14_io_macOut;
  wire       [7:0]    mac_5_15_io_passthrough;
  wire       [7:0]    mac_5_15_io_macOut;
  wire       [7:0]    mac_5_16_io_passthrough;
  wire       [7:0]    mac_5_16_io_macOut;
  wire       [7:0]    mac_5_17_io_passthrough;
  wire       [7:0]    mac_5_17_io_macOut;
  wire       [7:0]    mac_5_18_io_passthrough;
  wire       [7:0]    mac_5_18_io_macOut;
  wire       [7:0]    mac_5_19_io_passthrough;
  wire       [7:0]    mac_5_19_io_macOut;
  wire       [7:0]    mac_5_20_io_passthrough;
  wire       [7:0]    mac_5_20_io_macOut;
  wire       [7:0]    mac_5_21_io_passthrough;
  wire       [7:0]    mac_5_21_io_macOut;
  wire       [7:0]    mac_5_22_io_passthrough;
  wire       [7:0]    mac_5_22_io_macOut;
  wire       [7:0]    mac_5_23_io_passthrough;
  wire       [7:0]    mac_5_23_io_macOut;
  wire       [7:0]    mac_5_24_io_passthrough;
  wire       [7:0]    mac_5_24_io_macOut;
  wire       [7:0]    mac_5_25_io_passthrough;
  wire       [7:0]    mac_5_25_io_macOut;
  wire       [7:0]    mac_5_26_io_passthrough;
  wire       [7:0]    mac_5_26_io_macOut;
  wire       [7:0]    mac_5_27_io_passthrough;
  wire       [7:0]    mac_5_27_io_macOut;
  wire       [7:0]    mac_5_28_io_passthrough;
  wire       [7:0]    mac_5_28_io_macOut;
  wire       [7:0]    mac_5_29_io_passthrough;
  wire       [7:0]    mac_5_29_io_macOut;
  wire       [7:0]    mac_5_30_io_passthrough;
  wire       [7:0]    mac_5_30_io_macOut;
  wire       [7:0]    mac_5_31_io_passthrough;
  wire       [7:0]    mac_5_31_io_macOut;
  wire       [7:0]    mac_6_0_io_passthrough;
  wire       [7:0]    mac_6_0_io_macOut;
  wire       [7:0]    mac_6_1_io_passthrough;
  wire       [7:0]    mac_6_1_io_macOut;
  wire       [7:0]    mac_6_2_io_passthrough;
  wire       [7:0]    mac_6_2_io_macOut;
  wire       [7:0]    mac_6_3_io_passthrough;
  wire       [7:0]    mac_6_3_io_macOut;
  wire       [7:0]    mac_6_4_io_passthrough;
  wire       [7:0]    mac_6_4_io_macOut;
  wire       [7:0]    mac_6_5_io_passthrough;
  wire       [7:0]    mac_6_5_io_macOut;
  wire       [7:0]    mac_6_6_io_passthrough;
  wire       [7:0]    mac_6_6_io_macOut;
  wire       [7:0]    mac_6_7_io_passthrough;
  wire       [7:0]    mac_6_7_io_macOut;
  wire       [7:0]    mac_6_8_io_passthrough;
  wire       [7:0]    mac_6_8_io_macOut;
  wire       [7:0]    mac_6_9_io_passthrough;
  wire       [7:0]    mac_6_9_io_macOut;
  wire       [7:0]    mac_6_10_io_passthrough;
  wire       [7:0]    mac_6_10_io_macOut;
  wire       [7:0]    mac_6_11_io_passthrough;
  wire       [7:0]    mac_6_11_io_macOut;
  wire       [7:0]    mac_6_12_io_passthrough;
  wire       [7:0]    mac_6_12_io_macOut;
  wire       [7:0]    mac_6_13_io_passthrough;
  wire       [7:0]    mac_6_13_io_macOut;
  wire       [7:0]    mac_6_14_io_passthrough;
  wire       [7:0]    mac_6_14_io_macOut;
  wire       [7:0]    mac_6_15_io_passthrough;
  wire       [7:0]    mac_6_15_io_macOut;
  wire       [7:0]    mac_6_16_io_passthrough;
  wire       [7:0]    mac_6_16_io_macOut;
  wire       [7:0]    mac_6_17_io_passthrough;
  wire       [7:0]    mac_6_17_io_macOut;
  wire       [7:0]    mac_6_18_io_passthrough;
  wire       [7:0]    mac_6_18_io_macOut;
  wire       [7:0]    mac_6_19_io_passthrough;
  wire       [7:0]    mac_6_19_io_macOut;
  wire       [7:0]    mac_6_20_io_passthrough;
  wire       [7:0]    mac_6_20_io_macOut;
  wire       [7:0]    mac_6_21_io_passthrough;
  wire       [7:0]    mac_6_21_io_macOut;
  wire       [7:0]    mac_6_22_io_passthrough;
  wire       [7:0]    mac_6_22_io_macOut;
  wire       [7:0]    mac_6_23_io_passthrough;
  wire       [7:0]    mac_6_23_io_macOut;
  wire       [7:0]    mac_6_24_io_passthrough;
  wire       [7:0]    mac_6_24_io_macOut;
  wire       [7:0]    mac_6_25_io_passthrough;
  wire       [7:0]    mac_6_25_io_macOut;
  wire       [7:0]    mac_6_26_io_passthrough;
  wire       [7:0]    mac_6_26_io_macOut;
  wire       [7:0]    mac_6_27_io_passthrough;
  wire       [7:0]    mac_6_27_io_macOut;
  wire       [7:0]    mac_6_28_io_passthrough;
  wire       [7:0]    mac_6_28_io_macOut;
  wire       [7:0]    mac_6_29_io_passthrough;
  wire       [7:0]    mac_6_29_io_macOut;
  wire       [7:0]    mac_6_30_io_passthrough;
  wire       [7:0]    mac_6_30_io_macOut;
  wire       [7:0]    mac_6_31_io_passthrough;
  wire       [7:0]    mac_6_31_io_macOut;
  wire       [7:0]    mac_7_0_io_passthrough;
  wire       [7:0]    mac_7_0_io_macOut;
  wire       [7:0]    mac_7_1_io_passthrough;
  wire       [7:0]    mac_7_1_io_macOut;
  wire       [7:0]    mac_7_2_io_passthrough;
  wire       [7:0]    mac_7_2_io_macOut;
  wire       [7:0]    mac_7_3_io_passthrough;
  wire       [7:0]    mac_7_3_io_macOut;
  wire       [7:0]    mac_7_4_io_passthrough;
  wire       [7:0]    mac_7_4_io_macOut;
  wire       [7:0]    mac_7_5_io_passthrough;
  wire       [7:0]    mac_7_5_io_macOut;
  wire       [7:0]    mac_7_6_io_passthrough;
  wire       [7:0]    mac_7_6_io_macOut;
  wire       [7:0]    mac_7_7_io_passthrough;
  wire       [7:0]    mac_7_7_io_macOut;
  wire       [7:0]    mac_7_8_io_passthrough;
  wire       [7:0]    mac_7_8_io_macOut;
  wire       [7:0]    mac_7_9_io_passthrough;
  wire       [7:0]    mac_7_9_io_macOut;
  wire       [7:0]    mac_7_10_io_passthrough;
  wire       [7:0]    mac_7_10_io_macOut;
  wire       [7:0]    mac_7_11_io_passthrough;
  wire       [7:0]    mac_7_11_io_macOut;
  wire       [7:0]    mac_7_12_io_passthrough;
  wire       [7:0]    mac_7_12_io_macOut;
  wire       [7:0]    mac_7_13_io_passthrough;
  wire       [7:0]    mac_7_13_io_macOut;
  wire       [7:0]    mac_7_14_io_passthrough;
  wire       [7:0]    mac_7_14_io_macOut;
  wire       [7:0]    mac_7_15_io_passthrough;
  wire       [7:0]    mac_7_15_io_macOut;
  wire       [7:0]    mac_7_16_io_passthrough;
  wire       [7:0]    mac_7_16_io_macOut;
  wire       [7:0]    mac_7_17_io_passthrough;
  wire       [7:0]    mac_7_17_io_macOut;
  wire       [7:0]    mac_7_18_io_passthrough;
  wire       [7:0]    mac_7_18_io_macOut;
  wire       [7:0]    mac_7_19_io_passthrough;
  wire       [7:0]    mac_7_19_io_macOut;
  wire       [7:0]    mac_7_20_io_passthrough;
  wire       [7:0]    mac_7_20_io_macOut;
  wire       [7:0]    mac_7_21_io_passthrough;
  wire       [7:0]    mac_7_21_io_macOut;
  wire       [7:0]    mac_7_22_io_passthrough;
  wire       [7:0]    mac_7_22_io_macOut;
  wire       [7:0]    mac_7_23_io_passthrough;
  wire       [7:0]    mac_7_23_io_macOut;
  wire       [7:0]    mac_7_24_io_passthrough;
  wire       [7:0]    mac_7_24_io_macOut;
  wire       [7:0]    mac_7_25_io_passthrough;
  wire       [7:0]    mac_7_25_io_macOut;
  wire       [7:0]    mac_7_26_io_passthrough;
  wire       [7:0]    mac_7_26_io_macOut;
  wire       [7:0]    mac_7_27_io_passthrough;
  wire       [7:0]    mac_7_27_io_macOut;
  wire       [7:0]    mac_7_28_io_passthrough;
  wire       [7:0]    mac_7_28_io_macOut;
  wire       [7:0]    mac_7_29_io_passthrough;
  wire       [7:0]    mac_7_29_io_macOut;
  wire       [7:0]    mac_7_30_io_passthrough;
  wire       [7:0]    mac_7_30_io_macOut;
  wire       [7:0]    mac_7_31_io_passthrough;
  wire       [7:0]    mac_7_31_io_macOut;
  wire       [7:0]    mac_8_0_io_passthrough;
  wire       [7:0]    mac_8_0_io_macOut;
  wire       [7:0]    mac_8_1_io_passthrough;
  wire       [7:0]    mac_8_1_io_macOut;
  wire       [7:0]    mac_8_2_io_passthrough;
  wire       [7:0]    mac_8_2_io_macOut;
  wire       [7:0]    mac_8_3_io_passthrough;
  wire       [7:0]    mac_8_3_io_macOut;
  wire       [7:0]    mac_8_4_io_passthrough;
  wire       [7:0]    mac_8_4_io_macOut;
  wire       [7:0]    mac_8_5_io_passthrough;
  wire       [7:0]    mac_8_5_io_macOut;
  wire       [7:0]    mac_8_6_io_passthrough;
  wire       [7:0]    mac_8_6_io_macOut;
  wire       [7:0]    mac_8_7_io_passthrough;
  wire       [7:0]    mac_8_7_io_macOut;
  wire       [7:0]    mac_8_8_io_passthrough;
  wire       [7:0]    mac_8_8_io_macOut;
  wire       [7:0]    mac_8_9_io_passthrough;
  wire       [7:0]    mac_8_9_io_macOut;
  wire       [7:0]    mac_8_10_io_passthrough;
  wire       [7:0]    mac_8_10_io_macOut;
  wire       [7:0]    mac_8_11_io_passthrough;
  wire       [7:0]    mac_8_11_io_macOut;
  wire       [7:0]    mac_8_12_io_passthrough;
  wire       [7:0]    mac_8_12_io_macOut;
  wire       [7:0]    mac_8_13_io_passthrough;
  wire       [7:0]    mac_8_13_io_macOut;
  wire       [7:0]    mac_8_14_io_passthrough;
  wire       [7:0]    mac_8_14_io_macOut;
  wire       [7:0]    mac_8_15_io_passthrough;
  wire       [7:0]    mac_8_15_io_macOut;
  wire       [7:0]    mac_8_16_io_passthrough;
  wire       [7:0]    mac_8_16_io_macOut;
  wire       [7:0]    mac_8_17_io_passthrough;
  wire       [7:0]    mac_8_17_io_macOut;
  wire       [7:0]    mac_8_18_io_passthrough;
  wire       [7:0]    mac_8_18_io_macOut;
  wire       [7:0]    mac_8_19_io_passthrough;
  wire       [7:0]    mac_8_19_io_macOut;
  wire       [7:0]    mac_8_20_io_passthrough;
  wire       [7:0]    mac_8_20_io_macOut;
  wire       [7:0]    mac_8_21_io_passthrough;
  wire       [7:0]    mac_8_21_io_macOut;
  wire       [7:0]    mac_8_22_io_passthrough;
  wire       [7:0]    mac_8_22_io_macOut;
  wire       [7:0]    mac_8_23_io_passthrough;
  wire       [7:0]    mac_8_23_io_macOut;
  wire       [7:0]    mac_8_24_io_passthrough;
  wire       [7:0]    mac_8_24_io_macOut;
  wire       [7:0]    mac_8_25_io_passthrough;
  wire       [7:0]    mac_8_25_io_macOut;
  wire       [7:0]    mac_8_26_io_passthrough;
  wire       [7:0]    mac_8_26_io_macOut;
  wire       [7:0]    mac_8_27_io_passthrough;
  wire       [7:0]    mac_8_27_io_macOut;
  wire       [7:0]    mac_8_28_io_passthrough;
  wire       [7:0]    mac_8_28_io_macOut;
  wire       [7:0]    mac_8_29_io_passthrough;
  wire       [7:0]    mac_8_29_io_macOut;
  wire       [7:0]    mac_8_30_io_passthrough;
  wire       [7:0]    mac_8_30_io_macOut;
  wire       [7:0]    mac_8_31_io_passthrough;
  wire       [7:0]    mac_8_31_io_macOut;
  wire       [7:0]    mac_9_0_io_passthrough;
  wire       [7:0]    mac_9_0_io_macOut;
  wire       [7:0]    mac_9_1_io_passthrough;
  wire       [7:0]    mac_9_1_io_macOut;
  wire       [7:0]    mac_9_2_io_passthrough;
  wire       [7:0]    mac_9_2_io_macOut;
  wire       [7:0]    mac_9_3_io_passthrough;
  wire       [7:0]    mac_9_3_io_macOut;
  wire       [7:0]    mac_9_4_io_passthrough;
  wire       [7:0]    mac_9_4_io_macOut;
  wire       [7:0]    mac_9_5_io_passthrough;
  wire       [7:0]    mac_9_5_io_macOut;
  wire       [7:0]    mac_9_6_io_passthrough;
  wire       [7:0]    mac_9_6_io_macOut;
  wire       [7:0]    mac_9_7_io_passthrough;
  wire       [7:0]    mac_9_7_io_macOut;
  wire       [7:0]    mac_9_8_io_passthrough;
  wire       [7:0]    mac_9_8_io_macOut;
  wire       [7:0]    mac_9_9_io_passthrough;
  wire       [7:0]    mac_9_9_io_macOut;
  wire       [7:0]    mac_9_10_io_passthrough;
  wire       [7:0]    mac_9_10_io_macOut;
  wire       [7:0]    mac_9_11_io_passthrough;
  wire       [7:0]    mac_9_11_io_macOut;
  wire       [7:0]    mac_9_12_io_passthrough;
  wire       [7:0]    mac_9_12_io_macOut;
  wire       [7:0]    mac_9_13_io_passthrough;
  wire       [7:0]    mac_9_13_io_macOut;
  wire       [7:0]    mac_9_14_io_passthrough;
  wire       [7:0]    mac_9_14_io_macOut;
  wire       [7:0]    mac_9_15_io_passthrough;
  wire       [7:0]    mac_9_15_io_macOut;
  wire       [7:0]    mac_9_16_io_passthrough;
  wire       [7:0]    mac_9_16_io_macOut;
  wire       [7:0]    mac_9_17_io_passthrough;
  wire       [7:0]    mac_9_17_io_macOut;
  wire       [7:0]    mac_9_18_io_passthrough;
  wire       [7:0]    mac_9_18_io_macOut;
  wire       [7:0]    mac_9_19_io_passthrough;
  wire       [7:0]    mac_9_19_io_macOut;
  wire       [7:0]    mac_9_20_io_passthrough;
  wire       [7:0]    mac_9_20_io_macOut;
  wire       [7:0]    mac_9_21_io_passthrough;
  wire       [7:0]    mac_9_21_io_macOut;
  wire       [7:0]    mac_9_22_io_passthrough;
  wire       [7:0]    mac_9_22_io_macOut;
  wire       [7:0]    mac_9_23_io_passthrough;
  wire       [7:0]    mac_9_23_io_macOut;
  wire       [7:0]    mac_9_24_io_passthrough;
  wire       [7:0]    mac_9_24_io_macOut;
  wire       [7:0]    mac_9_25_io_passthrough;
  wire       [7:0]    mac_9_25_io_macOut;
  wire       [7:0]    mac_9_26_io_passthrough;
  wire       [7:0]    mac_9_26_io_macOut;
  wire       [7:0]    mac_9_27_io_passthrough;
  wire       [7:0]    mac_9_27_io_macOut;
  wire       [7:0]    mac_9_28_io_passthrough;
  wire       [7:0]    mac_9_28_io_macOut;
  wire       [7:0]    mac_9_29_io_passthrough;
  wire       [7:0]    mac_9_29_io_macOut;
  wire       [7:0]    mac_9_30_io_passthrough;
  wire       [7:0]    mac_9_30_io_macOut;
  wire       [7:0]    mac_9_31_io_passthrough;
  wire       [7:0]    mac_9_31_io_macOut;
  wire       [7:0]    mac_10_0_io_passthrough;
  wire       [7:0]    mac_10_0_io_macOut;
  wire       [7:0]    mac_10_1_io_passthrough;
  wire       [7:0]    mac_10_1_io_macOut;
  wire       [7:0]    mac_10_2_io_passthrough;
  wire       [7:0]    mac_10_2_io_macOut;
  wire       [7:0]    mac_10_3_io_passthrough;
  wire       [7:0]    mac_10_3_io_macOut;
  wire       [7:0]    mac_10_4_io_passthrough;
  wire       [7:0]    mac_10_4_io_macOut;
  wire       [7:0]    mac_10_5_io_passthrough;
  wire       [7:0]    mac_10_5_io_macOut;
  wire       [7:0]    mac_10_6_io_passthrough;
  wire       [7:0]    mac_10_6_io_macOut;
  wire       [7:0]    mac_10_7_io_passthrough;
  wire       [7:0]    mac_10_7_io_macOut;
  wire       [7:0]    mac_10_8_io_passthrough;
  wire       [7:0]    mac_10_8_io_macOut;
  wire       [7:0]    mac_10_9_io_passthrough;
  wire       [7:0]    mac_10_9_io_macOut;
  wire       [7:0]    mac_10_10_io_passthrough;
  wire       [7:0]    mac_10_10_io_macOut;
  wire       [7:0]    mac_10_11_io_passthrough;
  wire       [7:0]    mac_10_11_io_macOut;
  wire       [7:0]    mac_10_12_io_passthrough;
  wire       [7:0]    mac_10_12_io_macOut;
  wire       [7:0]    mac_10_13_io_passthrough;
  wire       [7:0]    mac_10_13_io_macOut;
  wire       [7:0]    mac_10_14_io_passthrough;
  wire       [7:0]    mac_10_14_io_macOut;
  wire       [7:0]    mac_10_15_io_passthrough;
  wire       [7:0]    mac_10_15_io_macOut;
  wire       [7:0]    mac_10_16_io_passthrough;
  wire       [7:0]    mac_10_16_io_macOut;
  wire       [7:0]    mac_10_17_io_passthrough;
  wire       [7:0]    mac_10_17_io_macOut;
  wire       [7:0]    mac_10_18_io_passthrough;
  wire       [7:0]    mac_10_18_io_macOut;
  wire       [7:0]    mac_10_19_io_passthrough;
  wire       [7:0]    mac_10_19_io_macOut;
  wire       [7:0]    mac_10_20_io_passthrough;
  wire       [7:0]    mac_10_20_io_macOut;
  wire       [7:0]    mac_10_21_io_passthrough;
  wire       [7:0]    mac_10_21_io_macOut;
  wire       [7:0]    mac_10_22_io_passthrough;
  wire       [7:0]    mac_10_22_io_macOut;
  wire       [7:0]    mac_10_23_io_passthrough;
  wire       [7:0]    mac_10_23_io_macOut;
  wire       [7:0]    mac_10_24_io_passthrough;
  wire       [7:0]    mac_10_24_io_macOut;
  wire       [7:0]    mac_10_25_io_passthrough;
  wire       [7:0]    mac_10_25_io_macOut;
  wire       [7:0]    mac_10_26_io_passthrough;
  wire       [7:0]    mac_10_26_io_macOut;
  wire       [7:0]    mac_10_27_io_passthrough;
  wire       [7:0]    mac_10_27_io_macOut;
  wire       [7:0]    mac_10_28_io_passthrough;
  wire       [7:0]    mac_10_28_io_macOut;
  wire       [7:0]    mac_10_29_io_passthrough;
  wire       [7:0]    mac_10_29_io_macOut;
  wire       [7:0]    mac_10_30_io_passthrough;
  wire       [7:0]    mac_10_30_io_macOut;
  wire       [7:0]    mac_10_31_io_passthrough;
  wire       [7:0]    mac_10_31_io_macOut;
  wire       [7:0]    mac_11_0_io_passthrough;
  wire       [7:0]    mac_11_0_io_macOut;
  wire       [7:0]    mac_11_1_io_passthrough;
  wire       [7:0]    mac_11_1_io_macOut;
  wire       [7:0]    mac_11_2_io_passthrough;
  wire       [7:0]    mac_11_2_io_macOut;
  wire       [7:0]    mac_11_3_io_passthrough;
  wire       [7:0]    mac_11_3_io_macOut;
  wire       [7:0]    mac_11_4_io_passthrough;
  wire       [7:0]    mac_11_4_io_macOut;
  wire       [7:0]    mac_11_5_io_passthrough;
  wire       [7:0]    mac_11_5_io_macOut;
  wire       [7:0]    mac_11_6_io_passthrough;
  wire       [7:0]    mac_11_6_io_macOut;
  wire       [7:0]    mac_11_7_io_passthrough;
  wire       [7:0]    mac_11_7_io_macOut;
  wire       [7:0]    mac_11_8_io_passthrough;
  wire       [7:0]    mac_11_8_io_macOut;
  wire       [7:0]    mac_11_9_io_passthrough;
  wire       [7:0]    mac_11_9_io_macOut;
  wire       [7:0]    mac_11_10_io_passthrough;
  wire       [7:0]    mac_11_10_io_macOut;
  wire       [7:0]    mac_11_11_io_passthrough;
  wire       [7:0]    mac_11_11_io_macOut;
  wire       [7:0]    mac_11_12_io_passthrough;
  wire       [7:0]    mac_11_12_io_macOut;
  wire       [7:0]    mac_11_13_io_passthrough;
  wire       [7:0]    mac_11_13_io_macOut;
  wire       [7:0]    mac_11_14_io_passthrough;
  wire       [7:0]    mac_11_14_io_macOut;
  wire       [7:0]    mac_11_15_io_passthrough;
  wire       [7:0]    mac_11_15_io_macOut;
  wire       [7:0]    mac_11_16_io_passthrough;
  wire       [7:0]    mac_11_16_io_macOut;
  wire       [7:0]    mac_11_17_io_passthrough;
  wire       [7:0]    mac_11_17_io_macOut;
  wire       [7:0]    mac_11_18_io_passthrough;
  wire       [7:0]    mac_11_18_io_macOut;
  wire       [7:0]    mac_11_19_io_passthrough;
  wire       [7:0]    mac_11_19_io_macOut;
  wire       [7:0]    mac_11_20_io_passthrough;
  wire       [7:0]    mac_11_20_io_macOut;
  wire       [7:0]    mac_11_21_io_passthrough;
  wire       [7:0]    mac_11_21_io_macOut;
  wire       [7:0]    mac_11_22_io_passthrough;
  wire       [7:0]    mac_11_22_io_macOut;
  wire       [7:0]    mac_11_23_io_passthrough;
  wire       [7:0]    mac_11_23_io_macOut;
  wire       [7:0]    mac_11_24_io_passthrough;
  wire       [7:0]    mac_11_24_io_macOut;
  wire       [7:0]    mac_11_25_io_passthrough;
  wire       [7:0]    mac_11_25_io_macOut;
  wire       [7:0]    mac_11_26_io_passthrough;
  wire       [7:0]    mac_11_26_io_macOut;
  wire       [7:0]    mac_11_27_io_passthrough;
  wire       [7:0]    mac_11_27_io_macOut;
  wire       [7:0]    mac_11_28_io_passthrough;
  wire       [7:0]    mac_11_28_io_macOut;
  wire       [7:0]    mac_11_29_io_passthrough;
  wire       [7:0]    mac_11_29_io_macOut;
  wire       [7:0]    mac_11_30_io_passthrough;
  wire       [7:0]    mac_11_30_io_macOut;
  wire       [7:0]    mac_11_31_io_passthrough;
  wire       [7:0]    mac_11_31_io_macOut;
  wire       [7:0]    mac_12_0_io_passthrough;
  wire       [7:0]    mac_12_0_io_macOut;
  wire       [7:0]    mac_12_1_io_passthrough;
  wire       [7:0]    mac_12_1_io_macOut;
  wire       [7:0]    mac_12_2_io_passthrough;
  wire       [7:0]    mac_12_2_io_macOut;
  wire       [7:0]    mac_12_3_io_passthrough;
  wire       [7:0]    mac_12_3_io_macOut;
  wire       [7:0]    mac_12_4_io_passthrough;
  wire       [7:0]    mac_12_4_io_macOut;
  wire       [7:0]    mac_12_5_io_passthrough;
  wire       [7:0]    mac_12_5_io_macOut;
  wire       [7:0]    mac_12_6_io_passthrough;
  wire       [7:0]    mac_12_6_io_macOut;
  wire       [7:0]    mac_12_7_io_passthrough;
  wire       [7:0]    mac_12_7_io_macOut;
  wire       [7:0]    mac_12_8_io_passthrough;
  wire       [7:0]    mac_12_8_io_macOut;
  wire       [7:0]    mac_12_9_io_passthrough;
  wire       [7:0]    mac_12_9_io_macOut;
  wire       [7:0]    mac_12_10_io_passthrough;
  wire       [7:0]    mac_12_10_io_macOut;
  wire       [7:0]    mac_12_11_io_passthrough;
  wire       [7:0]    mac_12_11_io_macOut;
  wire       [7:0]    mac_12_12_io_passthrough;
  wire       [7:0]    mac_12_12_io_macOut;
  wire       [7:0]    mac_12_13_io_passthrough;
  wire       [7:0]    mac_12_13_io_macOut;
  wire       [7:0]    mac_12_14_io_passthrough;
  wire       [7:0]    mac_12_14_io_macOut;
  wire       [7:0]    mac_12_15_io_passthrough;
  wire       [7:0]    mac_12_15_io_macOut;
  wire       [7:0]    mac_12_16_io_passthrough;
  wire       [7:0]    mac_12_16_io_macOut;
  wire       [7:0]    mac_12_17_io_passthrough;
  wire       [7:0]    mac_12_17_io_macOut;
  wire       [7:0]    mac_12_18_io_passthrough;
  wire       [7:0]    mac_12_18_io_macOut;
  wire       [7:0]    mac_12_19_io_passthrough;
  wire       [7:0]    mac_12_19_io_macOut;
  wire       [7:0]    mac_12_20_io_passthrough;
  wire       [7:0]    mac_12_20_io_macOut;
  wire       [7:0]    mac_12_21_io_passthrough;
  wire       [7:0]    mac_12_21_io_macOut;
  wire       [7:0]    mac_12_22_io_passthrough;
  wire       [7:0]    mac_12_22_io_macOut;
  wire       [7:0]    mac_12_23_io_passthrough;
  wire       [7:0]    mac_12_23_io_macOut;
  wire       [7:0]    mac_12_24_io_passthrough;
  wire       [7:0]    mac_12_24_io_macOut;
  wire       [7:0]    mac_12_25_io_passthrough;
  wire       [7:0]    mac_12_25_io_macOut;
  wire       [7:0]    mac_12_26_io_passthrough;
  wire       [7:0]    mac_12_26_io_macOut;
  wire       [7:0]    mac_12_27_io_passthrough;
  wire       [7:0]    mac_12_27_io_macOut;
  wire       [7:0]    mac_12_28_io_passthrough;
  wire       [7:0]    mac_12_28_io_macOut;
  wire       [7:0]    mac_12_29_io_passthrough;
  wire       [7:0]    mac_12_29_io_macOut;
  wire       [7:0]    mac_12_30_io_passthrough;
  wire       [7:0]    mac_12_30_io_macOut;
  wire       [7:0]    mac_12_31_io_passthrough;
  wire       [7:0]    mac_12_31_io_macOut;
  wire       [7:0]    mac_13_0_io_passthrough;
  wire       [7:0]    mac_13_0_io_macOut;
  wire       [7:0]    mac_13_1_io_passthrough;
  wire       [7:0]    mac_13_1_io_macOut;
  wire       [7:0]    mac_13_2_io_passthrough;
  wire       [7:0]    mac_13_2_io_macOut;
  wire       [7:0]    mac_13_3_io_passthrough;
  wire       [7:0]    mac_13_3_io_macOut;
  wire       [7:0]    mac_13_4_io_passthrough;
  wire       [7:0]    mac_13_4_io_macOut;
  wire       [7:0]    mac_13_5_io_passthrough;
  wire       [7:0]    mac_13_5_io_macOut;
  wire       [7:0]    mac_13_6_io_passthrough;
  wire       [7:0]    mac_13_6_io_macOut;
  wire       [7:0]    mac_13_7_io_passthrough;
  wire       [7:0]    mac_13_7_io_macOut;
  wire       [7:0]    mac_13_8_io_passthrough;
  wire       [7:0]    mac_13_8_io_macOut;
  wire       [7:0]    mac_13_9_io_passthrough;
  wire       [7:0]    mac_13_9_io_macOut;
  wire       [7:0]    mac_13_10_io_passthrough;
  wire       [7:0]    mac_13_10_io_macOut;
  wire       [7:0]    mac_13_11_io_passthrough;
  wire       [7:0]    mac_13_11_io_macOut;
  wire       [7:0]    mac_13_12_io_passthrough;
  wire       [7:0]    mac_13_12_io_macOut;
  wire       [7:0]    mac_13_13_io_passthrough;
  wire       [7:0]    mac_13_13_io_macOut;
  wire       [7:0]    mac_13_14_io_passthrough;
  wire       [7:0]    mac_13_14_io_macOut;
  wire       [7:0]    mac_13_15_io_passthrough;
  wire       [7:0]    mac_13_15_io_macOut;
  wire       [7:0]    mac_13_16_io_passthrough;
  wire       [7:0]    mac_13_16_io_macOut;
  wire       [7:0]    mac_13_17_io_passthrough;
  wire       [7:0]    mac_13_17_io_macOut;
  wire       [7:0]    mac_13_18_io_passthrough;
  wire       [7:0]    mac_13_18_io_macOut;
  wire       [7:0]    mac_13_19_io_passthrough;
  wire       [7:0]    mac_13_19_io_macOut;
  wire       [7:0]    mac_13_20_io_passthrough;
  wire       [7:0]    mac_13_20_io_macOut;
  wire       [7:0]    mac_13_21_io_passthrough;
  wire       [7:0]    mac_13_21_io_macOut;
  wire       [7:0]    mac_13_22_io_passthrough;
  wire       [7:0]    mac_13_22_io_macOut;
  wire       [7:0]    mac_13_23_io_passthrough;
  wire       [7:0]    mac_13_23_io_macOut;
  wire       [7:0]    mac_13_24_io_passthrough;
  wire       [7:0]    mac_13_24_io_macOut;
  wire       [7:0]    mac_13_25_io_passthrough;
  wire       [7:0]    mac_13_25_io_macOut;
  wire       [7:0]    mac_13_26_io_passthrough;
  wire       [7:0]    mac_13_26_io_macOut;
  wire       [7:0]    mac_13_27_io_passthrough;
  wire       [7:0]    mac_13_27_io_macOut;
  wire       [7:0]    mac_13_28_io_passthrough;
  wire       [7:0]    mac_13_28_io_macOut;
  wire       [7:0]    mac_13_29_io_passthrough;
  wire       [7:0]    mac_13_29_io_macOut;
  wire       [7:0]    mac_13_30_io_passthrough;
  wire       [7:0]    mac_13_30_io_macOut;
  wire       [7:0]    mac_13_31_io_passthrough;
  wire       [7:0]    mac_13_31_io_macOut;
  wire       [7:0]    mac_14_0_io_passthrough;
  wire       [7:0]    mac_14_0_io_macOut;
  wire       [7:0]    mac_14_1_io_passthrough;
  wire       [7:0]    mac_14_1_io_macOut;
  wire       [7:0]    mac_14_2_io_passthrough;
  wire       [7:0]    mac_14_2_io_macOut;
  wire       [7:0]    mac_14_3_io_passthrough;
  wire       [7:0]    mac_14_3_io_macOut;
  wire       [7:0]    mac_14_4_io_passthrough;
  wire       [7:0]    mac_14_4_io_macOut;
  wire       [7:0]    mac_14_5_io_passthrough;
  wire       [7:0]    mac_14_5_io_macOut;
  wire       [7:0]    mac_14_6_io_passthrough;
  wire       [7:0]    mac_14_6_io_macOut;
  wire       [7:0]    mac_14_7_io_passthrough;
  wire       [7:0]    mac_14_7_io_macOut;
  wire       [7:0]    mac_14_8_io_passthrough;
  wire       [7:0]    mac_14_8_io_macOut;
  wire       [7:0]    mac_14_9_io_passthrough;
  wire       [7:0]    mac_14_9_io_macOut;
  wire       [7:0]    mac_14_10_io_passthrough;
  wire       [7:0]    mac_14_10_io_macOut;
  wire       [7:0]    mac_14_11_io_passthrough;
  wire       [7:0]    mac_14_11_io_macOut;
  wire       [7:0]    mac_14_12_io_passthrough;
  wire       [7:0]    mac_14_12_io_macOut;
  wire       [7:0]    mac_14_13_io_passthrough;
  wire       [7:0]    mac_14_13_io_macOut;
  wire       [7:0]    mac_14_14_io_passthrough;
  wire       [7:0]    mac_14_14_io_macOut;
  wire       [7:0]    mac_14_15_io_passthrough;
  wire       [7:0]    mac_14_15_io_macOut;
  wire       [7:0]    mac_14_16_io_passthrough;
  wire       [7:0]    mac_14_16_io_macOut;
  wire       [7:0]    mac_14_17_io_passthrough;
  wire       [7:0]    mac_14_17_io_macOut;
  wire       [7:0]    mac_14_18_io_passthrough;
  wire       [7:0]    mac_14_18_io_macOut;
  wire       [7:0]    mac_14_19_io_passthrough;
  wire       [7:0]    mac_14_19_io_macOut;
  wire       [7:0]    mac_14_20_io_passthrough;
  wire       [7:0]    mac_14_20_io_macOut;
  wire       [7:0]    mac_14_21_io_passthrough;
  wire       [7:0]    mac_14_21_io_macOut;
  wire       [7:0]    mac_14_22_io_passthrough;
  wire       [7:0]    mac_14_22_io_macOut;
  wire       [7:0]    mac_14_23_io_passthrough;
  wire       [7:0]    mac_14_23_io_macOut;
  wire       [7:0]    mac_14_24_io_passthrough;
  wire       [7:0]    mac_14_24_io_macOut;
  wire       [7:0]    mac_14_25_io_passthrough;
  wire       [7:0]    mac_14_25_io_macOut;
  wire       [7:0]    mac_14_26_io_passthrough;
  wire       [7:0]    mac_14_26_io_macOut;
  wire       [7:0]    mac_14_27_io_passthrough;
  wire       [7:0]    mac_14_27_io_macOut;
  wire       [7:0]    mac_14_28_io_passthrough;
  wire       [7:0]    mac_14_28_io_macOut;
  wire       [7:0]    mac_14_29_io_passthrough;
  wire       [7:0]    mac_14_29_io_macOut;
  wire       [7:0]    mac_14_30_io_passthrough;
  wire       [7:0]    mac_14_30_io_macOut;
  wire       [7:0]    mac_14_31_io_passthrough;
  wire       [7:0]    mac_14_31_io_macOut;
  wire       [7:0]    mac_15_0_io_passthrough;
  wire       [7:0]    mac_15_0_io_macOut;
  wire       [7:0]    mac_15_1_io_passthrough;
  wire       [7:0]    mac_15_1_io_macOut;
  wire       [7:0]    mac_15_2_io_passthrough;
  wire       [7:0]    mac_15_2_io_macOut;
  wire       [7:0]    mac_15_3_io_passthrough;
  wire       [7:0]    mac_15_3_io_macOut;
  wire       [7:0]    mac_15_4_io_passthrough;
  wire       [7:0]    mac_15_4_io_macOut;
  wire       [7:0]    mac_15_5_io_passthrough;
  wire       [7:0]    mac_15_5_io_macOut;
  wire       [7:0]    mac_15_6_io_passthrough;
  wire       [7:0]    mac_15_6_io_macOut;
  wire       [7:0]    mac_15_7_io_passthrough;
  wire       [7:0]    mac_15_7_io_macOut;
  wire       [7:0]    mac_15_8_io_passthrough;
  wire       [7:0]    mac_15_8_io_macOut;
  wire       [7:0]    mac_15_9_io_passthrough;
  wire       [7:0]    mac_15_9_io_macOut;
  wire       [7:0]    mac_15_10_io_passthrough;
  wire       [7:0]    mac_15_10_io_macOut;
  wire       [7:0]    mac_15_11_io_passthrough;
  wire       [7:0]    mac_15_11_io_macOut;
  wire       [7:0]    mac_15_12_io_passthrough;
  wire       [7:0]    mac_15_12_io_macOut;
  wire       [7:0]    mac_15_13_io_passthrough;
  wire       [7:0]    mac_15_13_io_macOut;
  wire       [7:0]    mac_15_14_io_passthrough;
  wire       [7:0]    mac_15_14_io_macOut;
  wire       [7:0]    mac_15_15_io_passthrough;
  wire       [7:0]    mac_15_15_io_macOut;
  wire       [7:0]    mac_15_16_io_passthrough;
  wire       [7:0]    mac_15_16_io_macOut;
  wire       [7:0]    mac_15_17_io_passthrough;
  wire       [7:0]    mac_15_17_io_macOut;
  wire       [7:0]    mac_15_18_io_passthrough;
  wire       [7:0]    mac_15_18_io_macOut;
  wire       [7:0]    mac_15_19_io_passthrough;
  wire       [7:0]    mac_15_19_io_macOut;
  wire       [7:0]    mac_15_20_io_passthrough;
  wire       [7:0]    mac_15_20_io_macOut;
  wire       [7:0]    mac_15_21_io_passthrough;
  wire       [7:0]    mac_15_21_io_macOut;
  wire       [7:0]    mac_15_22_io_passthrough;
  wire       [7:0]    mac_15_22_io_macOut;
  wire       [7:0]    mac_15_23_io_passthrough;
  wire       [7:0]    mac_15_23_io_macOut;
  wire       [7:0]    mac_15_24_io_passthrough;
  wire       [7:0]    mac_15_24_io_macOut;
  wire       [7:0]    mac_15_25_io_passthrough;
  wire       [7:0]    mac_15_25_io_macOut;
  wire       [7:0]    mac_15_26_io_passthrough;
  wire       [7:0]    mac_15_26_io_macOut;
  wire       [7:0]    mac_15_27_io_passthrough;
  wire       [7:0]    mac_15_27_io_macOut;
  wire       [7:0]    mac_15_28_io_passthrough;
  wire       [7:0]    mac_15_28_io_macOut;
  wire       [7:0]    mac_15_29_io_passthrough;
  wire       [7:0]    mac_15_29_io_macOut;
  wire       [7:0]    mac_15_30_io_passthrough;
  wire       [7:0]    mac_15_30_io_macOut;
  wire       [7:0]    mac_15_31_io_passthrough;
  wire       [7:0]    mac_15_31_io_macOut;
  wire       [7:0]    mac_16_0_io_passthrough;
  wire       [7:0]    mac_16_0_io_macOut;
  wire       [7:0]    mac_16_1_io_passthrough;
  wire       [7:0]    mac_16_1_io_macOut;
  wire       [7:0]    mac_16_2_io_passthrough;
  wire       [7:0]    mac_16_2_io_macOut;
  wire       [7:0]    mac_16_3_io_passthrough;
  wire       [7:0]    mac_16_3_io_macOut;
  wire       [7:0]    mac_16_4_io_passthrough;
  wire       [7:0]    mac_16_4_io_macOut;
  wire       [7:0]    mac_16_5_io_passthrough;
  wire       [7:0]    mac_16_5_io_macOut;
  wire       [7:0]    mac_16_6_io_passthrough;
  wire       [7:0]    mac_16_6_io_macOut;
  wire       [7:0]    mac_16_7_io_passthrough;
  wire       [7:0]    mac_16_7_io_macOut;
  wire       [7:0]    mac_16_8_io_passthrough;
  wire       [7:0]    mac_16_8_io_macOut;
  wire       [7:0]    mac_16_9_io_passthrough;
  wire       [7:0]    mac_16_9_io_macOut;
  wire       [7:0]    mac_16_10_io_passthrough;
  wire       [7:0]    mac_16_10_io_macOut;
  wire       [7:0]    mac_16_11_io_passthrough;
  wire       [7:0]    mac_16_11_io_macOut;
  wire       [7:0]    mac_16_12_io_passthrough;
  wire       [7:0]    mac_16_12_io_macOut;
  wire       [7:0]    mac_16_13_io_passthrough;
  wire       [7:0]    mac_16_13_io_macOut;
  wire       [7:0]    mac_16_14_io_passthrough;
  wire       [7:0]    mac_16_14_io_macOut;
  wire       [7:0]    mac_16_15_io_passthrough;
  wire       [7:0]    mac_16_15_io_macOut;
  wire       [7:0]    mac_16_16_io_passthrough;
  wire       [7:0]    mac_16_16_io_macOut;
  wire       [7:0]    mac_16_17_io_passthrough;
  wire       [7:0]    mac_16_17_io_macOut;
  wire       [7:0]    mac_16_18_io_passthrough;
  wire       [7:0]    mac_16_18_io_macOut;
  wire       [7:0]    mac_16_19_io_passthrough;
  wire       [7:0]    mac_16_19_io_macOut;
  wire       [7:0]    mac_16_20_io_passthrough;
  wire       [7:0]    mac_16_20_io_macOut;
  wire       [7:0]    mac_16_21_io_passthrough;
  wire       [7:0]    mac_16_21_io_macOut;
  wire       [7:0]    mac_16_22_io_passthrough;
  wire       [7:0]    mac_16_22_io_macOut;
  wire       [7:0]    mac_16_23_io_passthrough;
  wire       [7:0]    mac_16_23_io_macOut;
  wire       [7:0]    mac_16_24_io_passthrough;
  wire       [7:0]    mac_16_24_io_macOut;
  wire       [7:0]    mac_16_25_io_passthrough;
  wire       [7:0]    mac_16_25_io_macOut;
  wire       [7:0]    mac_16_26_io_passthrough;
  wire       [7:0]    mac_16_26_io_macOut;
  wire       [7:0]    mac_16_27_io_passthrough;
  wire       [7:0]    mac_16_27_io_macOut;
  wire       [7:0]    mac_16_28_io_passthrough;
  wire       [7:0]    mac_16_28_io_macOut;
  wire       [7:0]    mac_16_29_io_passthrough;
  wire       [7:0]    mac_16_29_io_macOut;
  wire       [7:0]    mac_16_30_io_passthrough;
  wire       [7:0]    mac_16_30_io_macOut;
  wire       [7:0]    mac_16_31_io_passthrough;
  wire       [7:0]    mac_16_31_io_macOut;
  wire       [7:0]    mac_17_0_io_passthrough;
  wire       [7:0]    mac_17_0_io_macOut;
  wire       [7:0]    mac_17_1_io_passthrough;
  wire       [7:0]    mac_17_1_io_macOut;
  wire       [7:0]    mac_17_2_io_passthrough;
  wire       [7:0]    mac_17_2_io_macOut;
  wire       [7:0]    mac_17_3_io_passthrough;
  wire       [7:0]    mac_17_3_io_macOut;
  wire       [7:0]    mac_17_4_io_passthrough;
  wire       [7:0]    mac_17_4_io_macOut;
  wire       [7:0]    mac_17_5_io_passthrough;
  wire       [7:0]    mac_17_5_io_macOut;
  wire       [7:0]    mac_17_6_io_passthrough;
  wire       [7:0]    mac_17_6_io_macOut;
  wire       [7:0]    mac_17_7_io_passthrough;
  wire       [7:0]    mac_17_7_io_macOut;
  wire       [7:0]    mac_17_8_io_passthrough;
  wire       [7:0]    mac_17_8_io_macOut;
  wire       [7:0]    mac_17_9_io_passthrough;
  wire       [7:0]    mac_17_9_io_macOut;
  wire       [7:0]    mac_17_10_io_passthrough;
  wire       [7:0]    mac_17_10_io_macOut;
  wire       [7:0]    mac_17_11_io_passthrough;
  wire       [7:0]    mac_17_11_io_macOut;
  wire       [7:0]    mac_17_12_io_passthrough;
  wire       [7:0]    mac_17_12_io_macOut;
  wire       [7:0]    mac_17_13_io_passthrough;
  wire       [7:0]    mac_17_13_io_macOut;
  wire       [7:0]    mac_17_14_io_passthrough;
  wire       [7:0]    mac_17_14_io_macOut;
  wire       [7:0]    mac_17_15_io_passthrough;
  wire       [7:0]    mac_17_15_io_macOut;
  wire       [7:0]    mac_17_16_io_passthrough;
  wire       [7:0]    mac_17_16_io_macOut;
  wire       [7:0]    mac_17_17_io_passthrough;
  wire       [7:0]    mac_17_17_io_macOut;
  wire       [7:0]    mac_17_18_io_passthrough;
  wire       [7:0]    mac_17_18_io_macOut;
  wire       [7:0]    mac_17_19_io_passthrough;
  wire       [7:0]    mac_17_19_io_macOut;
  wire       [7:0]    mac_17_20_io_passthrough;
  wire       [7:0]    mac_17_20_io_macOut;
  wire       [7:0]    mac_17_21_io_passthrough;
  wire       [7:0]    mac_17_21_io_macOut;
  wire       [7:0]    mac_17_22_io_passthrough;
  wire       [7:0]    mac_17_22_io_macOut;
  wire       [7:0]    mac_17_23_io_passthrough;
  wire       [7:0]    mac_17_23_io_macOut;
  wire       [7:0]    mac_17_24_io_passthrough;
  wire       [7:0]    mac_17_24_io_macOut;
  wire       [7:0]    mac_17_25_io_passthrough;
  wire       [7:0]    mac_17_25_io_macOut;
  wire       [7:0]    mac_17_26_io_passthrough;
  wire       [7:0]    mac_17_26_io_macOut;
  wire       [7:0]    mac_17_27_io_passthrough;
  wire       [7:0]    mac_17_27_io_macOut;
  wire       [7:0]    mac_17_28_io_passthrough;
  wire       [7:0]    mac_17_28_io_macOut;
  wire       [7:0]    mac_17_29_io_passthrough;
  wire       [7:0]    mac_17_29_io_macOut;
  wire       [7:0]    mac_17_30_io_passthrough;
  wire       [7:0]    mac_17_30_io_macOut;
  wire       [7:0]    mac_17_31_io_passthrough;
  wire       [7:0]    mac_17_31_io_macOut;
  wire       [7:0]    mac_18_0_io_passthrough;
  wire       [7:0]    mac_18_0_io_macOut;
  wire       [7:0]    mac_18_1_io_passthrough;
  wire       [7:0]    mac_18_1_io_macOut;
  wire       [7:0]    mac_18_2_io_passthrough;
  wire       [7:0]    mac_18_2_io_macOut;
  wire       [7:0]    mac_18_3_io_passthrough;
  wire       [7:0]    mac_18_3_io_macOut;
  wire       [7:0]    mac_18_4_io_passthrough;
  wire       [7:0]    mac_18_4_io_macOut;
  wire       [7:0]    mac_18_5_io_passthrough;
  wire       [7:0]    mac_18_5_io_macOut;
  wire       [7:0]    mac_18_6_io_passthrough;
  wire       [7:0]    mac_18_6_io_macOut;
  wire       [7:0]    mac_18_7_io_passthrough;
  wire       [7:0]    mac_18_7_io_macOut;
  wire       [7:0]    mac_18_8_io_passthrough;
  wire       [7:0]    mac_18_8_io_macOut;
  wire       [7:0]    mac_18_9_io_passthrough;
  wire       [7:0]    mac_18_9_io_macOut;
  wire       [7:0]    mac_18_10_io_passthrough;
  wire       [7:0]    mac_18_10_io_macOut;
  wire       [7:0]    mac_18_11_io_passthrough;
  wire       [7:0]    mac_18_11_io_macOut;
  wire       [7:0]    mac_18_12_io_passthrough;
  wire       [7:0]    mac_18_12_io_macOut;
  wire       [7:0]    mac_18_13_io_passthrough;
  wire       [7:0]    mac_18_13_io_macOut;
  wire       [7:0]    mac_18_14_io_passthrough;
  wire       [7:0]    mac_18_14_io_macOut;
  wire       [7:0]    mac_18_15_io_passthrough;
  wire       [7:0]    mac_18_15_io_macOut;
  wire       [7:0]    mac_18_16_io_passthrough;
  wire       [7:0]    mac_18_16_io_macOut;
  wire       [7:0]    mac_18_17_io_passthrough;
  wire       [7:0]    mac_18_17_io_macOut;
  wire       [7:0]    mac_18_18_io_passthrough;
  wire       [7:0]    mac_18_18_io_macOut;
  wire       [7:0]    mac_18_19_io_passthrough;
  wire       [7:0]    mac_18_19_io_macOut;
  wire       [7:0]    mac_18_20_io_passthrough;
  wire       [7:0]    mac_18_20_io_macOut;
  wire       [7:0]    mac_18_21_io_passthrough;
  wire       [7:0]    mac_18_21_io_macOut;
  wire       [7:0]    mac_18_22_io_passthrough;
  wire       [7:0]    mac_18_22_io_macOut;
  wire       [7:0]    mac_18_23_io_passthrough;
  wire       [7:0]    mac_18_23_io_macOut;
  wire       [7:0]    mac_18_24_io_passthrough;
  wire       [7:0]    mac_18_24_io_macOut;
  wire       [7:0]    mac_18_25_io_passthrough;
  wire       [7:0]    mac_18_25_io_macOut;
  wire       [7:0]    mac_18_26_io_passthrough;
  wire       [7:0]    mac_18_26_io_macOut;
  wire       [7:0]    mac_18_27_io_passthrough;
  wire       [7:0]    mac_18_27_io_macOut;
  wire       [7:0]    mac_18_28_io_passthrough;
  wire       [7:0]    mac_18_28_io_macOut;
  wire       [7:0]    mac_18_29_io_passthrough;
  wire       [7:0]    mac_18_29_io_macOut;
  wire       [7:0]    mac_18_30_io_passthrough;
  wire       [7:0]    mac_18_30_io_macOut;
  wire       [7:0]    mac_18_31_io_passthrough;
  wire       [7:0]    mac_18_31_io_macOut;
  wire       [7:0]    mac_19_0_io_passthrough;
  wire       [7:0]    mac_19_0_io_macOut;
  wire       [7:0]    mac_19_1_io_passthrough;
  wire       [7:0]    mac_19_1_io_macOut;
  wire       [7:0]    mac_19_2_io_passthrough;
  wire       [7:0]    mac_19_2_io_macOut;
  wire       [7:0]    mac_19_3_io_passthrough;
  wire       [7:0]    mac_19_3_io_macOut;
  wire       [7:0]    mac_19_4_io_passthrough;
  wire       [7:0]    mac_19_4_io_macOut;
  wire       [7:0]    mac_19_5_io_passthrough;
  wire       [7:0]    mac_19_5_io_macOut;
  wire       [7:0]    mac_19_6_io_passthrough;
  wire       [7:0]    mac_19_6_io_macOut;
  wire       [7:0]    mac_19_7_io_passthrough;
  wire       [7:0]    mac_19_7_io_macOut;
  wire       [7:0]    mac_19_8_io_passthrough;
  wire       [7:0]    mac_19_8_io_macOut;
  wire       [7:0]    mac_19_9_io_passthrough;
  wire       [7:0]    mac_19_9_io_macOut;
  wire       [7:0]    mac_19_10_io_passthrough;
  wire       [7:0]    mac_19_10_io_macOut;
  wire       [7:0]    mac_19_11_io_passthrough;
  wire       [7:0]    mac_19_11_io_macOut;
  wire       [7:0]    mac_19_12_io_passthrough;
  wire       [7:0]    mac_19_12_io_macOut;
  wire       [7:0]    mac_19_13_io_passthrough;
  wire       [7:0]    mac_19_13_io_macOut;
  wire       [7:0]    mac_19_14_io_passthrough;
  wire       [7:0]    mac_19_14_io_macOut;
  wire       [7:0]    mac_19_15_io_passthrough;
  wire       [7:0]    mac_19_15_io_macOut;
  wire       [7:0]    mac_19_16_io_passthrough;
  wire       [7:0]    mac_19_16_io_macOut;
  wire       [7:0]    mac_19_17_io_passthrough;
  wire       [7:0]    mac_19_17_io_macOut;
  wire       [7:0]    mac_19_18_io_passthrough;
  wire       [7:0]    mac_19_18_io_macOut;
  wire       [7:0]    mac_19_19_io_passthrough;
  wire       [7:0]    mac_19_19_io_macOut;
  wire       [7:0]    mac_19_20_io_passthrough;
  wire       [7:0]    mac_19_20_io_macOut;
  wire       [7:0]    mac_19_21_io_passthrough;
  wire       [7:0]    mac_19_21_io_macOut;
  wire       [7:0]    mac_19_22_io_passthrough;
  wire       [7:0]    mac_19_22_io_macOut;
  wire       [7:0]    mac_19_23_io_passthrough;
  wire       [7:0]    mac_19_23_io_macOut;
  wire       [7:0]    mac_19_24_io_passthrough;
  wire       [7:0]    mac_19_24_io_macOut;
  wire       [7:0]    mac_19_25_io_passthrough;
  wire       [7:0]    mac_19_25_io_macOut;
  wire       [7:0]    mac_19_26_io_passthrough;
  wire       [7:0]    mac_19_26_io_macOut;
  wire       [7:0]    mac_19_27_io_passthrough;
  wire       [7:0]    mac_19_27_io_macOut;
  wire       [7:0]    mac_19_28_io_passthrough;
  wire       [7:0]    mac_19_28_io_macOut;
  wire       [7:0]    mac_19_29_io_passthrough;
  wire       [7:0]    mac_19_29_io_macOut;
  wire       [7:0]    mac_19_30_io_passthrough;
  wire       [7:0]    mac_19_30_io_macOut;
  wire       [7:0]    mac_19_31_io_passthrough;
  wire       [7:0]    mac_19_31_io_macOut;
  wire       [7:0]    mac_20_0_io_passthrough;
  wire       [7:0]    mac_20_0_io_macOut;
  wire       [7:0]    mac_20_1_io_passthrough;
  wire       [7:0]    mac_20_1_io_macOut;
  wire       [7:0]    mac_20_2_io_passthrough;
  wire       [7:0]    mac_20_2_io_macOut;
  wire       [7:0]    mac_20_3_io_passthrough;
  wire       [7:0]    mac_20_3_io_macOut;
  wire       [7:0]    mac_20_4_io_passthrough;
  wire       [7:0]    mac_20_4_io_macOut;
  wire       [7:0]    mac_20_5_io_passthrough;
  wire       [7:0]    mac_20_5_io_macOut;
  wire       [7:0]    mac_20_6_io_passthrough;
  wire       [7:0]    mac_20_6_io_macOut;
  wire       [7:0]    mac_20_7_io_passthrough;
  wire       [7:0]    mac_20_7_io_macOut;
  wire       [7:0]    mac_20_8_io_passthrough;
  wire       [7:0]    mac_20_8_io_macOut;
  wire       [7:0]    mac_20_9_io_passthrough;
  wire       [7:0]    mac_20_9_io_macOut;
  wire       [7:0]    mac_20_10_io_passthrough;
  wire       [7:0]    mac_20_10_io_macOut;
  wire       [7:0]    mac_20_11_io_passthrough;
  wire       [7:0]    mac_20_11_io_macOut;
  wire       [7:0]    mac_20_12_io_passthrough;
  wire       [7:0]    mac_20_12_io_macOut;
  wire       [7:0]    mac_20_13_io_passthrough;
  wire       [7:0]    mac_20_13_io_macOut;
  wire       [7:0]    mac_20_14_io_passthrough;
  wire       [7:0]    mac_20_14_io_macOut;
  wire       [7:0]    mac_20_15_io_passthrough;
  wire       [7:0]    mac_20_15_io_macOut;
  wire       [7:0]    mac_20_16_io_passthrough;
  wire       [7:0]    mac_20_16_io_macOut;
  wire       [7:0]    mac_20_17_io_passthrough;
  wire       [7:0]    mac_20_17_io_macOut;
  wire       [7:0]    mac_20_18_io_passthrough;
  wire       [7:0]    mac_20_18_io_macOut;
  wire       [7:0]    mac_20_19_io_passthrough;
  wire       [7:0]    mac_20_19_io_macOut;
  wire       [7:0]    mac_20_20_io_passthrough;
  wire       [7:0]    mac_20_20_io_macOut;
  wire       [7:0]    mac_20_21_io_passthrough;
  wire       [7:0]    mac_20_21_io_macOut;
  wire       [7:0]    mac_20_22_io_passthrough;
  wire       [7:0]    mac_20_22_io_macOut;
  wire       [7:0]    mac_20_23_io_passthrough;
  wire       [7:0]    mac_20_23_io_macOut;
  wire       [7:0]    mac_20_24_io_passthrough;
  wire       [7:0]    mac_20_24_io_macOut;
  wire       [7:0]    mac_20_25_io_passthrough;
  wire       [7:0]    mac_20_25_io_macOut;
  wire       [7:0]    mac_20_26_io_passthrough;
  wire       [7:0]    mac_20_26_io_macOut;
  wire       [7:0]    mac_20_27_io_passthrough;
  wire       [7:0]    mac_20_27_io_macOut;
  wire       [7:0]    mac_20_28_io_passthrough;
  wire       [7:0]    mac_20_28_io_macOut;
  wire       [7:0]    mac_20_29_io_passthrough;
  wire       [7:0]    mac_20_29_io_macOut;
  wire       [7:0]    mac_20_30_io_passthrough;
  wire       [7:0]    mac_20_30_io_macOut;
  wire       [7:0]    mac_20_31_io_passthrough;
  wire       [7:0]    mac_20_31_io_macOut;
  wire       [7:0]    mac_21_0_io_passthrough;
  wire       [7:0]    mac_21_0_io_macOut;
  wire       [7:0]    mac_21_1_io_passthrough;
  wire       [7:0]    mac_21_1_io_macOut;
  wire       [7:0]    mac_21_2_io_passthrough;
  wire       [7:0]    mac_21_2_io_macOut;
  wire       [7:0]    mac_21_3_io_passthrough;
  wire       [7:0]    mac_21_3_io_macOut;
  wire       [7:0]    mac_21_4_io_passthrough;
  wire       [7:0]    mac_21_4_io_macOut;
  wire       [7:0]    mac_21_5_io_passthrough;
  wire       [7:0]    mac_21_5_io_macOut;
  wire       [7:0]    mac_21_6_io_passthrough;
  wire       [7:0]    mac_21_6_io_macOut;
  wire       [7:0]    mac_21_7_io_passthrough;
  wire       [7:0]    mac_21_7_io_macOut;
  wire       [7:0]    mac_21_8_io_passthrough;
  wire       [7:0]    mac_21_8_io_macOut;
  wire       [7:0]    mac_21_9_io_passthrough;
  wire       [7:0]    mac_21_9_io_macOut;
  wire       [7:0]    mac_21_10_io_passthrough;
  wire       [7:0]    mac_21_10_io_macOut;
  wire       [7:0]    mac_21_11_io_passthrough;
  wire       [7:0]    mac_21_11_io_macOut;
  wire       [7:0]    mac_21_12_io_passthrough;
  wire       [7:0]    mac_21_12_io_macOut;
  wire       [7:0]    mac_21_13_io_passthrough;
  wire       [7:0]    mac_21_13_io_macOut;
  wire       [7:0]    mac_21_14_io_passthrough;
  wire       [7:0]    mac_21_14_io_macOut;
  wire       [7:0]    mac_21_15_io_passthrough;
  wire       [7:0]    mac_21_15_io_macOut;
  wire       [7:0]    mac_21_16_io_passthrough;
  wire       [7:0]    mac_21_16_io_macOut;
  wire       [7:0]    mac_21_17_io_passthrough;
  wire       [7:0]    mac_21_17_io_macOut;
  wire       [7:0]    mac_21_18_io_passthrough;
  wire       [7:0]    mac_21_18_io_macOut;
  wire       [7:0]    mac_21_19_io_passthrough;
  wire       [7:0]    mac_21_19_io_macOut;
  wire       [7:0]    mac_21_20_io_passthrough;
  wire       [7:0]    mac_21_20_io_macOut;
  wire       [7:0]    mac_21_21_io_passthrough;
  wire       [7:0]    mac_21_21_io_macOut;
  wire       [7:0]    mac_21_22_io_passthrough;
  wire       [7:0]    mac_21_22_io_macOut;
  wire       [7:0]    mac_21_23_io_passthrough;
  wire       [7:0]    mac_21_23_io_macOut;
  wire       [7:0]    mac_21_24_io_passthrough;
  wire       [7:0]    mac_21_24_io_macOut;
  wire       [7:0]    mac_21_25_io_passthrough;
  wire       [7:0]    mac_21_25_io_macOut;
  wire       [7:0]    mac_21_26_io_passthrough;
  wire       [7:0]    mac_21_26_io_macOut;
  wire       [7:0]    mac_21_27_io_passthrough;
  wire       [7:0]    mac_21_27_io_macOut;
  wire       [7:0]    mac_21_28_io_passthrough;
  wire       [7:0]    mac_21_28_io_macOut;
  wire       [7:0]    mac_21_29_io_passthrough;
  wire       [7:0]    mac_21_29_io_macOut;
  wire       [7:0]    mac_21_30_io_passthrough;
  wire       [7:0]    mac_21_30_io_macOut;
  wire       [7:0]    mac_21_31_io_passthrough;
  wire       [7:0]    mac_21_31_io_macOut;
  wire       [7:0]    mac_22_0_io_passthrough;
  wire       [7:0]    mac_22_0_io_macOut;
  wire       [7:0]    mac_22_1_io_passthrough;
  wire       [7:0]    mac_22_1_io_macOut;
  wire       [7:0]    mac_22_2_io_passthrough;
  wire       [7:0]    mac_22_2_io_macOut;
  wire       [7:0]    mac_22_3_io_passthrough;
  wire       [7:0]    mac_22_3_io_macOut;
  wire       [7:0]    mac_22_4_io_passthrough;
  wire       [7:0]    mac_22_4_io_macOut;
  wire       [7:0]    mac_22_5_io_passthrough;
  wire       [7:0]    mac_22_5_io_macOut;
  wire       [7:0]    mac_22_6_io_passthrough;
  wire       [7:0]    mac_22_6_io_macOut;
  wire       [7:0]    mac_22_7_io_passthrough;
  wire       [7:0]    mac_22_7_io_macOut;
  wire       [7:0]    mac_22_8_io_passthrough;
  wire       [7:0]    mac_22_8_io_macOut;
  wire       [7:0]    mac_22_9_io_passthrough;
  wire       [7:0]    mac_22_9_io_macOut;
  wire       [7:0]    mac_22_10_io_passthrough;
  wire       [7:0]    mac_22_10_io_macOut;
  wire       [7:0]    mac_22_11_io_passthrough;
  wire       [7:0]    mac_22_11_io_macOut;
  wire       [7:0]    mac_22_12_io_passthrough;
  wire       [7:0]    mac_22_12_io_macOut;
  wire       [7:0]    mac_22_13_io_passthrough;
  wire       [7:0]    mac_22_13_io_macOut;
  wire       [7:0]    mac_22_14_io_passthrough;
  wire       [7:0]    mac_22_14_io_macOut;
  wire       [7:0]    mac_22_15_io_passthrough;
  wire       [7:0]    mac_22_15_io_macOut;
  wire       [7:0]    mac_22_16_io_passthrough;
  wire       [7:0]    mac_22_16_io_macOut;
  wire       [7:0]    mac_22_17_io_passthrough;
  wire       [7:0]    mac_22_17_io_macOut;
  wire       [7:0]    mac_22_18_io_passthrough;
  wire       [7:0]    mac_22_18_io_macOut;
  wire       [7:0]    mac_22_19_io_passthrough;
  wire       [7:0]    mac_22_19_io_macOut;
  wire       [7:0]    mac_22_20_io_passthrough;
  wire       [7:0]    mac_22_20_io_macOut;
  wire       [7:0]    mac_22_21_io_passthrough;
  wire       [7:0]    mac_22_21_io_macOut;
  wire       [7:0]    mac_22_22_io_passthrough;
  wire       [7:0]    mac_22_22_io_macOut;
  wire       [7:0]    mac_22_23_io_passthrough;
  wire       [7:0]    mac_22_23_io_macOut;
  wire       [7:0]    mac_22_24_io_passthrough;
  wire       [7:0]    mac_22_24_io_macOut;
  wire       [7:0]    mac_22_25_io_passthrough;
  wire       [7:0]    mac_22_25_io_macOut;
  wire       [7:0]    mac_22_26_io_passthrough;
  wire       [7:0]    mac_22_26_io_macOut;
  wire       [7:0]    mac_22_27_io_passthrough;
  wire       [7:0]    mac_22_27_io_macOut;
  wire       [7:0]    mac_22_28_io_passthrough;
  wire       [7:0]    mac_22_28_io_macOut;
  wire       [7:0]    mac_22_29_io_passthrough;
  wire       [7:0]    mac_22_29_io_macOut;
  wire       [7:0]    mac_22_30_io_passthrough;
  wire       [7:0]    mac_22_30_io_macOut;
  wire       [7:0]    mac_22_31_io_passthrough;
  wire       [7:0]    mac_22_31_io_macOut;
  wire       [7:0]    mac_23_0_io_passthrough;
  wire       [7:0]    mac_23_0_io_macOut;
  wire       [7:0]    mac_23_1_io_passthrough;
  wire       [7:0]    mac_23_1_io_macOut;
  wire       [7:0]    mac_23_2_io_passthrough;
  wire       [7:0]    mac_23_2_io_macOut;
  wire       [7:0]    mac_23_3_io_passthrough;
  wire       [7:0]    mac_23_3_io_macOut;
  wire       [7:0]    mac_23_4_io_passthrough;
  wire       [7:0]    mac_23_4_io_macOut;
  wire       [7:0]    mac_23_5_io_passthrough;
  wire       [7:0]    mac_23_5_io_macOut;
  wire       [7:0]    mac_23_6_io_passthrough;
  wire       [7:0]    mac_23_6_io_macOut;
  wire       [7:0]    mac_23_7_io_passthrough;
  wire       [7:0]    mac_23_7_io_macOut;
  wire       [7:0]    mac_23_8_io_passthrough;
  wire       [7:0]    mac_23_8_io_macOut;
  wire       [7:0]    mac_23_9_io_passthrough;
  wire       [7:0]    mac_23_9_io_macOut;
  wire       [7:0]    mac_23_10_io_passthrough;
  wire       [7:0]    mac_23_10_io_macOut;
  wire       [7:0]    mac_23_11_io_passthrough;
  wire       [7:0]    mac_23_11_io_macOut;
  wire       [7:0]    mac_23_12_io_passthrough;
  wire       [7:0]    mac_23_12_io_macOut;
  wire       [7:0]    mac_23_13_io_passthrough;
  wire       [7:0]    mac_23_13_io_macOut;
  wire       [7:0]    mac_23_14_io_passthrough;
  wire       [7:0]    mac_23_14_io_macOut;
  wire       [7:0]    mac_23_15_io_passthrough;
  wire       [7:0]    mac_23_15_io_macOut;
  wire       [7:0]    mac_23_16_io_passthrough;
  wire       [7:0]    mac_23_16_io_macOut;
  wire       [7:0]    mac_23_17_io_passthrough;
  wire       [7:0]    mac_23_17_io_macOut;
  wire       [7:0]    mac_23_18_io_passthrough;
  wire       [7:0]    mac_23_18_io_macOut;
  wire       [7:0]    mac_23_19_io_passthrough;
  wire       [7:0]    mac_23_19_io_macOut;
  wire       [7:0]    mac_23_20_io_passthrough;
  wire       [7:0]    mac_23_20_io_macOut;
  wire       [7:0]    mac_23_21_io_passthrough;
  wire       [7:0]    mac_23_21_io_macOut;
  wire       [7:0]    mac_23_22_io_passthrough;
  wire       [7:0]    mac_23_22_io_macOut;
  wire       [7:0]    mac_23_23_io_passthrough;
  wire       [7:0]    mac_23_23_io_macOut;
  wire       [7:0]    mac_23_24_io_passthrough;
  wire       [7:0]    mac_23_24_io_macOut;
  wire       [7:0]    mac_23_25_io_passthrough;
  wire       [7:0]    mac_23_25_io_macOut;
  wire       [7:0]    mac_23_26_io_passthrough;
  wire       [7:0]    mac_23_26_io_macOut;
  wire       [7:0]    mac_23_27_io_passthrough;
  wire       [7:0]    mac_23_27_io_macOut;
  wire       [7:0]    mac_23_28_io_passthrough;
  wire       [7:0]    mac_23_28_io_macOut;
  wire       [7:0]    mac_23_29_io_passthrough;
  wire       [7:0]    mac_23_29_io_macOut;
  wire       [7:0]    mac_23_30_io_passthrough;
  wire       [7:0]    mac_23_30_io_macOut;
  wire       [7:0]    mac_23_31_io_passthrough;
  wire       [7:0]    mac_23_31_io_macOut;
  wire       [7:0]    mac_24_0_io_passthrough;
  wire       [7:0]    mac_24_0_io_macOut;
  wire       [7:0]    mac_24_1_io_passthrough;
  wire       [7:0]    mac_24_1_io_macOut;
  wire       [7:0]    mac_24_2_io_passthrough;
  wire       [7:0]    mac_24_2_io_macOut;
  wire       [7:0]    mac_24_3_io_passthrough;
  wire       [7:0]    mac_24_3_io_macOut;
  wire       [7:0]    mac_24_4_io_passthrough;
  wire       [7:0]    mac_24_4_io_macOut;
  wire       [7:0]    mac_24_5_io_passthrough;
  wire       [7:0]    mac_24_5_io_macOut;
  wire       [7:0]    mac_24_6_io_passthrough;
  wire       [7:0]    mac_24_6_io_macOut;
  wire       [7:0]    mac_24_7_io_passthrough;
  wire       [7:0]    mac_24_7_io_macOut;
  wire       [7:0]    mac_24_8_io_passthrough;
  wire       [7:0]    mac_24_8_io_macOut;
  wire       [7:0]    mac_24_9_io_passthrough;
  wire       [7:0]    mac_24_9_io_macOut;
  wire       [7:0]    mac_24_10_io_passthrough;
  wire       [7:0]    mac_24_10_io_macOut;
  wire       [7:0]    mac_24_11_io_passthrough;
  wire       [7:0]    mac_24_11_io_macOut;
  wire       [7:0]    mac_24_12_io_passthrough;
  wire       [7:0]    mac_24_12_io_macOut;
  wire       [7:0]    mac_24_13_io_passthrough;
  wire       [7:0]    mac_24_13_io_macOut;
  wire       [7:0]    mac_24_14_io_passthrough;
  wire       [7:0]    mac_24_14_io_macOut;
  wire       [7:0]    mac_24_15_io_passthrough;
  wire       [7:0]    mac_24_15_io_macOut;
  wire       [7:0]    mac_24_16_io_passthrough;
  wire       [7:0]    mac_24_16_io_macOut;
  wire       [7:0]    mac_24_17_io_passthrough;
  wire       [7:0]    mac_24_17_io_macOut;
  wire       [7:0]    mac_24_18_io_passthrough;
  wire       [7:0]    mac_24_18_io_macOut;
  wire       [7:0]    mac_24_19_io_passthrough;
  wire       [7:0]    mac_24_19_io_macOut;
  wire       [7:0]    mac_24_20_io_passthrough;
  wire       [7:0]    mac_24_20_io_macOut;
  wire       [7:0]    mac_24_21_io_passthrough;
  wire       [7:0]    mac_24_21_io_macOut;
  wire       [7:0]    mac_24_22_io_passthrough;
  wire       [7:0]    mac_24_22_io_macOut;
  wire       [7:0]    mac_24_23_io_passthrough;
  wire       [7:0]    mac_24_23_io_macOut;
  wire       [7:0]    mac_24_24_io_passthrough;
  wire       [7:0]    mac_24_24_io_macOut;
  wire       [7:0]    mac_24_25_io_passthrough;
  wire       [7:0]    mac_24_25_io_macOut;
  wire       [7:0]    mac_24_26_io_passthrough;
  wire       [7:0]    mac_24_26_io_macOut;
  wire       [7:0]    mac_24_27_io_passthrough;
  wire       [7:0]    mac_24_27_io_macOut;
  wire       [7:0]    mac_24_28_io_passthrough;
  wire       [7:0]    mac_24_28_io_macOut;
  wire       [7:0]    mac_24_29_io_passthrough;
  wire       [7:0]    mac_24_29_io_macOut;
  wire       [7:0]    mac_24_30_io_passthrough;
  wire       [7:0]    mac_24_30_io_macOut;
  wire       [7:0]    mac_24_31_io_passthrough;
  wire       [7:0]    mac_24_31_io_macOut;
  wire       [7:0]    mac_25_0_io_passthrough;
  wire       [7:0]    mac_25_0_io_macOut;
  wire       [7:0]    mac_25_1_io_passthrough;
  wire       [7:0]    mac_25_1_io_macOut;
  wire       [7:0]    mac_25_2_io_passthrough;
  wire       [7:0]    mac_25_2_io_macOut;
  wire       [7:0]    mac_25_3_io_passthrough;
  wire       [7:0]    mac_25_3_io_macOut;
  wire       [7:0]    mac_25_4_io_passthrough;
  wire       [7:0]    mac_25_4_io_macOut;
  wire       [7:0]    mac_25_5_io_passthrough;
  wire       [7:0]    mac_25_5_io_macOut;
  wire       [7:0]    mac_25_6_io_passthrough;
  wire       [7:0]    mac_25_6_io_macOut;
  wire       [7:0]    mac_25_7_io_passthrough;
  wire       [7:0]    mac_25_7_io_macOut;
  wire       [7:0]    mac_25_8_io_passthrough;
  wire       [7:0]    mac_25_8_io_macOut;
  wire       [7:0]    mac_25_9_io_passthrough;
  wire       [7:0]    mac_25_9_io_macOut;
  wire       [7:0]    mac_25_10_io_passthrough;
  wire       [7:0]    mac_25_10_io_macOut;
  wire       [7:0]    mac_25_11_io_passthrough;
  wire       [7:0]    mac_25_11_io_macOut;
  wire       [7:0]    mac_25_12_io_passthrough;
  wire       [7:0]    mac_25_12_io_macOut;
  wire       [7:0]    mac_25_13_io_passthrough;
  wire       [7:0]    mac_25_13_io_macOut;
  wire       [7:0]    mac_25_14_io_passthrough;
  wire       [7:0]    mac_25_14_io_macOut;
  wire       [7:0]    mac_25_15_io_passthrough;
  wire       [7:0]    mac_25_15_io_macOut;
  wire       [7:0]    mac_25_16_io_passthrough;
  wire       [7:0]    mac_25_16_io_macOut;
  wire       [7:0]    mac_25_17_io_passthrough;
  wire       [7:0]    mac_25_17_io_macOut;
  wire       [7:0]    mac_25_18_io_passthrough;
  wire       [7:0]    mac_25_18_io_macOut;
  wire       [7:0]    mac_25_19_io_passthrough;
  wire       [7:0]    mac_25_19_io_macOut;
  wire       [7:0]    mac_25_20_io_passthrough;
  wire       [7:0]    mac_25_20_io_macOut;
  wire       [7:0]    mac_25_21_io_passthrough;
  wire       [7:0]    mac_25_21_io_macOut;
  wire       [7:0]    mac_25_22_io_passthrough;
  wire       [7:0]    mac_25_22_io_macOut;
  wire       [7:0]    mac_25_23_io_passthrough;
  wire       [7:0]    mac_25_23_io_macOut;
  wire       [7:0]    mac_25_24_io_passthrough;
  wire       [7:0]    mac_25_24_io_macOut;
  wire       [7:0]    mac_25_25_io_passthrough;
  wire       [7:0]    mac_25_25_io_macOut;
  wire       [7:0]    mac_25_26_io_passthrough;
  wire       [7:0]    mac_25_26_io_macOut;
  wire       [7:0]    mac_25_27_io_passthrough;
  wire       [7:0]    mac_25_27_io_macOut;
  wire       [7:0]    mac_25_28_io_passthrough;
  wire       [7:0]    mac_25_28_io_macOut;
  wire       [7:0]    mac_25_29_io_passthrough;
  wire       [7:0]    mac_25_29_io_macOut;
  wire       [7:0]    mac_25_30_io_passthrough;
  wire       [7:0]    mac_25_30_io_macOut;
  wire       [7:0]    mac_25_31_io_passthrough;
  wire       [7:0]    mac_25_31_io_macOut;
  wire       [7:0]    mac_26_0_io_passthrough;
  wire       [7:0]    mac_26_0_io_macOut;
  wire       [7:0]    mac_26_1_io_passthrough;
  wire       [7:0]    mac_26_1_io_macOut;
  wire       [7:0]    mac_26_2_io_passthrough;
  wire       [7:0]    mac_26_2_io_macOut;
  wire       [7:0]    mac_26_3_io_passthrough;
  wire       [7:0]    mac_26_3_io_macOut;
  wire       [7:0]    mac_26_4_io_passthrough;
  wire       [7:0]    mac_26_4_io_macOut;
  wire       [7:0]    mac_26_5_io_passthrough;
  wire       [7:0]    mac_26_5_io_macOut;
  wire       [7:0]    mac_26_6_io_passthrough;
  wire       [7:0]    mac_26_6_io_macOut;
  wire       [7:0]    mac_26_7_io_passthrough;
  wire       [7:0]    mac_26_7_io_macOut;
  wire       [7:0]    mac_26_8_io_passthrough;
  wire       [7:0]    mac_26_8_io_macOut;
  wire       [7:0]    mac_26_9_io_passthrough;
  wire       [7:0]    mac_26_9_io_macOut;
  wire       [7:0]    mac_26_10_io_passthrough;
  wire       [7:0]    mac_26_10_io_macOut;
  wire       [7:0]    mac_26_11_io_passthrough;
  wire       [7:0]    mac_26_11_io_macOut;
  wire       [7:0]    mac_26_12_io_passthrough;
  wire       [7:0]    mac_26_12_io_macOut;
  wire       [7:0]    mac_26_13_io_passthrough;
  wire       [7:0]    mac_26_13_io_macOut;
  wire       [7:0]    mac_26_14_io_passthrough;
  wire       [7:0]    mac_26_14_io_macOut;
  wire       [7:0]    mac_26_15_io_passthrough;
  wire       [7:0]    mac_26_15_io_macOut;
  wire       [7:0]    mac_26_16_io_passthrough;
  wire       [7:0]    mac_26_16_io_macOut;
  wire       [7:0]    mac_26_17_io_passthrough;
  wire       [7:0]    mac_26_17_io_macOut;
  wire       [7:0]    mac_26_18_io_passthrough;
  wire       [7:0]    mac_26_18_io_macOut;
  wire       [7:0]    mac_26_19_io_passthrough;
  wire       [7:0]    mac_26_19_io_macOut;
  wire       [7:0]    mac_26_20_io_passthrough;
  wire       [7:0]    mac_26_20_io_macOut;
  wire       [7:0]    mac_26_21_io_passthrough;
  wire       [7:0]    mac_26_21_io_macOut;
  wire       [7:0]    mac_26_22_io_passthrough;
  wire       [7:0]    mac_26_22_io_macOut;
  wire       [7:0]    mac_26_23_io_passthrough;
  wire       [7:0]    mac_26_23_io_macOut;
  wire       [7:0]    mac_26_24_io_passthrough;
  wire       [7:0]    mac_26_24_io_macOut;
  wire       [7:0]    mac_26_25_io_passthrough;
  wire       [7:0]    mac_26_25_io_macOut;
  wire       [7:0]    mac_26_26_io_passthrough;
  wire       [7:0]    mac_26_26_io_macOut;
  wire       [7:0]    mac_26_27_io_passthrough;
  wire       [7:0]    mac_26_27_io_macOut;
  wire       [7:0]    mac_26_28_io_passthrough;
  wire       [7:0]    mac_26_28_io_macOut;
  wire       [7:0]    mac_26_29_io_passthrough;
  wire       [7:0]    mac_26_29_io_macOut;
  wire       [7:0]    mac_26_30_io_passthrough;
  wire       [7:0]    mac_26_30_io_macOut;
  wire       [7:0]    mac_26_31_io_passthrough;
  wire       [7:0]    mac_26_31_io_macOut;
  wire       [7:0]    mac_27_0_io_passthrough;
  wire       [7:0]    mac_27_0_io_macOut;
  wire       [7:0]    mac_27_1_io_passthrough;
  wire       [7:0]    mac_27_1_io_macOut;
  wire       [7:0]    mac_27_2_io_passthrough;
  wire       [7:0]    mac_27_2_io_macOut;
  wire       [7:0]    mac_27_3_io_passthrough;
  wire       [7:0]    mac_27_3_io_macOut;
  wire       [7:0]    mac_27_4_io_passthrough;
  wire       [7:0]    mac_27_4_io_macOut;
  wire       [7:0]    mac_27_5_io_passthrough;
  wire       [7:0]    mac_27_5_io_macOut;
  wire       [7:0]    mac_27_6_io_passthrough;
  wire       [7:0]    mac_27_6_io_macOut;
  wire       [7:0]    mac_27_7_io_passthrough;
  wire       [7:0]    mac_27_7_io_macOut;
  wire       [7:0]    mac_27_8_io_passthrough;
  wire       [7:0]    mac_27_8_io_macOut;
  wire       [7:0]    mac_27_9_io_passthrough;
  wire       [7:0]    mac_27_9_io_macOut;
  wire       [7:0]    mac_27_10_io_passthrough;
  wire       [7:0]    mac_27_10_io_macOut;
  wire       [7:0]    mac_27_11_io_passthrough;
  wire       [7:0]    mac_27_11_io_macOut;
  wire       [7:0]    mac_27_12_io_passthrough;
  wire       [7:0]    mac_27_12_io_macOut;
  wire       [7:0]    mac_27_13_io_passthrough;
  wire       [7:0]    mac_27_13_io_macOut;
  wire       [7:0]    mac_27_14_io_passthrough;
  wire       [7:0]    mac_27_14_io_macOut;
  wire       [7:0]    mac_27_15_io_passthrough;
  wire       [7:0]    mac_27_15_io_macOut;
  wire       [7:0]    mac_27_16_io_passthrough;
  wire       [7:0]    mac_27_16_io_macOut;
  wire       [7:0]    mac_27_17_io_passthrough;
  wire       [7:0]    mac_27_17_io_macOut;
  wire       [7:0]    mac_27_18_io_passthrough;
  wire       [7:0]    mac_27_18_io_macOut;
  wire       [7:0]    mac_27_19_io_passthrough;
  wire       [7:0]    mac_27_19_io_macOut;
  wire       [7:0]    mac_27_20_io_passthrough;
  wire       [7:0]    mac_27_20_io_macOut;
  wire       [7:0]    mac_27_21_io_passthrough;
  wire       [7:0]    mac_27_21_io_macOut;
  wire       [7:0]    mac_27_22_io_passthrough;
  wire       [7:0]    mac_27_22_io_macOut;
  wire       [7:0]    mac_27_23_io_passthrough;
  wire       [7:0]    mac_27_23_io_macOut;
  wire       [7:0]    mac_27_24_io_passthrough;
  wire       [7:0]    mac_27_24_io_macOut;
  wire       [7:0]    mac_27_25_io_passthrough;
  wire       [7:0]    mac_27_25_io_macOut;
  wire       [7:0]    mac_27_26_io_passthrough;
  wire       [7:0]    mac_27_26_io_macOut;
  wire       [7:0]    mac_27_27_io_passthrough;
  wire       [7:0]    mac_27_27_io_macOut;
  wire       [7:0]    mac_27_28_io_passthrough;
  wire       [7:0]    mac_27_28_io_macOut;
  wire       [7:0]    mac_27_29_io_passthrough;
  wire       [7:0]    mac_27_29_io_macOut;
  wire       [7:0]    mac_27_30_io_passthrough;
  wire       [7:0]    mac_27_30_io_macOut;
  wire       [7:0]    mac_27_31_io_passthrough;
  wire       [7:0]    mac_27_31_io_macOut;
  wire       [7:0]    mac_28_0_io_passthrough;
  wire       [7:0]    mac_28_0_io_macOut;
  wire       [7:0]    mac_28_1_io_passthrough;
  wire       [7:0]    mac_28_1_io_macOut;
  wire       [7:0]    mac_28_2_io_passthrough;
  wire       [7:0]    mac_28_2_io_macOut;
  wire       [7:0]    mac_28_3_io_passthrough;
  wire       [7:0]    mac_28_3_io_macOut;
  wire       [7:0]    mac_28_4_io_passthrough;
  wire       [7:0]    mac_28_4_io_macOut;
  wire       [7:0]    mac_28_5_io_passthrough;
  wire       [7:0]    mac_28_5_io_macOut;
  wire       [7:0]    mac_28_6_io_passthrough;
  wire       [7:0]    mac_28_6_io_macOut;
  wire       [7:0]    mac_28_7_io_passthrough;
  wire       [7:0]    mac_28_7_io_macOut;
  wire       [7:0]    mac_28_8_io_passthrough;
  wire       [7:0]    mac_28_8_io_macOut;
  wire       [7:0]    mac_28_9_io_passthrough;
  wire       [7:0]    mac_28_9_io_macOut;
  wire       [7:0]    mac_28_10_io_passthrough;
  wire       [7:0]    mac_28_10_io_macOut;
  wire       [7:0]    mac_28_11_io_passthrough;
  wire       [7:0]    mac_28_11_io_macOut;
  wire       [7:0]    mac_28_12_io_passthrough;
  wire       [7:0]    mac_28_12_io_macOut;
  wire       [7:0]    mac_28_13_io_passthrough;
  wire       [7:0]    mac_28_13_io_macOut;
  wire       [7:0]    mac_28_14_io_passthrough;
  wire       [7:0]    mac_28_14_io_macOut;
  wire       [7:0]    mac_28_15_io_passthrough;
  wire       [7:0]    mac_28_15_io_macOut;
  wire       [7:0]    mac_28_16_io_passthrough;
  wire       [7:0]    mac_28_16_io_macOut;
  wire       [7:0]    mac_28_17_io_passthrough;
  wire       [7:0]    mac_28_17_io_macOut;
  wire       [7:0]    mac_28_18_io_passthrough;
  wire       [7:0]    mac_28_18_io_macOut;
  wire       [7:0]    mac_28_19_io_passthrough;
  wire       [7:0]    mac_28_19_io_macOut;
  wire       [7:0]    mac_28_20_io_passthrough;
  wire       [7:0]    mac_28_20_io_macOut;
  wire       [7:0]    mac_28_21_io_passthrough;
  wire       [7:0]    mac_28_21_io_macOut;
  wire       [7:0]    mac_28_22_io_passthrough;
  wire       [7:0]    mac_28_22_io_macOut;
  wire       [7:0]    mac_28_23_io_passthrough;
  wire       [7:0]    mac_28_23_io_macOut;
  wire       [7:0]    mac_28_24_io_passthrough;
  wire       [7:0]    mac_28_24_io_macOut;
  wire       [7:0]    mac_28_25_io_passthrough;
  wire       [7:0]    mac_28_25_io_macOut;
  wire       [7:0]    mac_28_26_io_passthrough;
  wire       [7:0]    mac_28_26_io_macOut;
  wire       [7:0]    mac_28_27_io_passthrough;
  wire       [7:0]    mac_28_27_io_macOut;
  wire       [7:0]    mac_28_28_io_passthrough;
  wire       [7:0]    mac_28_28_io_macOut;
  wire       [7:0]    mac_28_29_io_passthrough;
  wire       [7:0]    mac_28_29_io_macOut;
  wire       [7:0]    mac_28_30_io_passthrough;
  wire       [7:0]    mac_28_30_io_macOut;
  wire       [7:0]    mac_28_31_io_passthrough;
  wire       [7:0]    mac_28_31_io_macOut;
  wire       [7:0]    mac_29_0_io_passthrough;
  wire       [7:0]    mac_29_0_io_macOut;
  wire       [7:0]    mac_29_1_io_passthrough;
  wire       [7:0]    mac_29_1_io_macOut;
  wire       [7:0]    mac_29_2_io_passthrough;
  wire       [7:0]    mac_29_2_io_macOut;
  wire       [7:0]    mac_29_3_io_passthrough;
  wire       [7:0]    mac_29_3_io_macOut;
  wire       [7:0]    mac_29_4_io_passthrough;
  wire       [7:0]    mac_29_4_io_macOut;
  wire       [7:0]    mac_29_5_io_passthrough;
  wire       [7:0]    mac_29_5_io_macOut;
  wire       [7:0]    mac_29_6_io_passthrough;
  wire       [7:0]    mac_29_6_io_macOut;
  wire       [7:0]    mac_29_7_io_passthrough;
  wire       [7:0]    mac_29_7_io_macOut;
  wire       [7:0]    mac_29_8_io_passthrough;
  wire       [7:0]    mac_29_8_io_macOut;
  wire       [7:0]    mac_29_9_io_passthrough;
  wire       [7:0]    mac_29_9_io_macOut;
  wire       [7:0]    mac_29_10_io_passthrough;
  wire       [7:0]    mac_29_10_io_macOut;
  wire       [7:0]    mac_29_11_io_passthrough;
  wire       [7:0]    mac_29_11_io_macOut;
  wire       [7:0]    mac_29_12_io_passthrough;
  wire       [7:0]    mac_29_12_io_macOut;
  wire       [7:0]    mac_29_13_io_passthrough;
  wire       [7:0]    mac_29_13_io_macOut;
  wire       [7:0]    mac_29_14_io_passthrough;
  wire       [7:0]    mac_29_14_io_macOut;
  wire       [7:0]    mac_29_15_io_passthrough;
  wire       [7:0]    mac_29_15_io_macOut;
  wire       [7:0]    mac_29_16_io_passthrough;
  wire       [7:0]    mac_29_16_io_macOut;
  wire       [7:0]    mac_29_17_io_passthrough;
  wire       [7:0]    mac_29_17_io_macOut;
  wire       [7:0]    mac_29_18_io_passthrough;
  wire       [7:0]    mac_29_18_io_macOut;
  wire       [7:0]    mac_29_19_io_passthrough;
  wire       [7:0]    mac_29_19_io_macOut;
  wire       [7:0]    mac_29_20_io_passthrough;
  wire       [7:0]    mac_29_20_io_macOut;
  wire       [7:0]    mac_29_21_io_passthrough;
  wire       [7:0]    mac_29_21_io_macOut;
  wire       [7:0]    mac_29_22_io_passthrough;
  wire       [7:0]    mac_29_22_io_macOut;
  wire       [7:0]    mac_29_23_io_passthrough;
  wire       [7:0]    mac_29_23_io_macOut;
  wire       [7:0]    mac_29_24_io_passthrough;
  wire       [7:0]    mac_29_24_io_macOut;
  wire       [7:0]    mac_29_25_io_passthrough;
  wire       [7:0]    mac_29_25_io_macOut;
  wire       [7:0]    mac_29_26_io_passthrough;
  wire       [7:0]    mac_29_26_io_macOut;
  wire       [7:0]    mac_29_27_io_passthrough;
  wire       [7:0]    mac_29_27_io_macOut;
  wire       [7:0]    mac_29_28_io_passthrough;
  wire       [7:0]    mac_29_28_io_macOut;
  wire       [7:0]    mac_29_29_io_passthrough;
  wire       [7:0]    mac_29_29_io_macOut;
  wire       [7:0]    mac_29_30_io_passthrough;
  wire       [7:0]    mac_29_30_io_macOut;
  wire       [7:0]    mac_29_31_io_passthrough;
  wire       [7:0]    mac_29_31_io_macOut;
  wire       [7:0]    mac_30_0_io_passthrough;
  wire       [7:0]    mac_30_0_io_macOut;
  wire       [7:0]    mac_30_1_io_passthrough;
  wire       [7:0]    mac_30_1_io_macOut;
  wire       [7:0]    mac_30_2_io_passthrough;
  wire       [7:0]    mac_30_2_io_macOut;
  wire       [7:0]    mac_30_3_io_passthrough;
  wire       [7:0]    mac_30_3_io_macOut;
  wire       [7:0]    mac_30_4_io_passthrough;
  wire       [7:0]    mac_30_4_io_macOut;
  wire       [7:0]    mac_30_5_io_passthrough;
  wire       [7:0]    mac_30_5_io_macOut;
  wire       [7:0]    mac_30_6_io_passthrough;
  wire       [7:0]    mac_30_6_io_macOut;
  wire       [7:0]    mac_30_7_io_passthrough;
  wire       [7:0]    mac_30_7_io_macOut;
  wire       [7:0]    mac_30_8_io_passthrough;
  wire       [7:0]    mac_30_8_io_macOut;
  wire       [7:0]    mac_30_9_io_passthrough;
  wire       [7:0]    mac_30_9_io_macOut;
  wire       [7:0]    mac_30_10_io_passthrough;
  wire       [7:0]    mac_30_10_io_macOut;
  wire       [7:0]    mac_30_11_io_passthrough;
  wire       [7:0]    mac_30_11_io_macOut;
  wire       [7:0]    mac_30_12_io_passthrough;
  wire       [7:0]    mac_30_12_io_macOut;
  wire       [7:0]    mac_30_13_io_passthrough;
  wire       [7:0]    mac_30_13_io_macOut;
  wire       [7:0]    mac_30_14_io_passthrough;
  wire       [7:0]    mac_30_14_io_macOut;
  wire       [7:0]    mac_30_15_io_passthrough;
  wire       [7:0]    mac_30_15_io_macOut;
  wire       [7:0]    mac_30_16_io_passthrough;
  wire       [7:0]    mac_30_16_io_macOut;
  wire       [7:0]    mac_30_17_io_passthrough;
  wire       [7:0]    mac_30_17_io_macOut;
  wire       [7:0]    mac_30_18_io_passthrough;
  wire       [7:0]    mac_30_18_io_macOut;
  wire       [7:0]    mac_30_19_io_passthrough;
  wire       [7:0]    mac_30_19_io_macOut;
  wire       [7:0]    mac_30_20_io_passthrough;
  wire       [7:0]    mac_30_20_io_macOut;
  wire       [7:0]    mac_30_21_io_passthrough;
  wire       [7:0]    mac_30_21_io_macOut;
  wire       [7:0]    mac_30_22_io_passthrough;
  wire       [7:0]    mac_30_22_io_macOut;
  wire       [7:0]    mac_30_23_io_passthrough;
  wire       [7:0]    mac_30_23_io_macOut;
  wire       [7:0]    mac_30_24_io_passthrough;
  wire       [7:0]    mac_30_24_io_macOut;
  wire       [7:0]    mac_30_25_io_passthrough;
  wire       [7:0]    mac_30_25_io_macOut;
  wire       [7:0]    mac_30_26_io_passthrough;
  wire       [7:0]    mac_30_26_io_macOut;
  wire       [7:0]    mac_30_27_io_passthrough;
  wire       [7:0]    mac_30_27_io_macOut;
  wire       [7:0]    mac_30_28_io_passthrough;
  wire       [7:0]    mac_30_28_io_macOut;
  wire       [7:0]    mac_30_29_io_passthrough;
  wire       [7:0]    mac_30_29_io_macOut;
  wire       [7:0]    mac_30_30_io_passthrough;
  wire       [7:0]    mac_30_30_io_macOut;
  wire       [7:0]    mac_30_31_io_passthrough;
  wire       [7:0]    mac_30_31_io_macOut;
  wire       [7:0]    mac_31_0_io_passthrough;
  wire       [7:0]    mac_31_0_io_macOut;
  wire       [7:0]    mac_31_1_io_passthrough;
  wire       [7:0]    mac_31_1_io_macOut;
  wire       [7:0]    mac_31_2_io_passthrough;
  wire       [7:0]    mac_31_2_io_macOut;
  wire       [7:0]    mac_31_3_io_passthrough;
  wire       [7:0]    mac_31_3_io_macOut;
  wire       [7:0]    mac_31_4_io_passthrough;
  wire       [7:0]    mac_31_4_io_macOut;
  wire       [7:0]    mac_31_5_io_passthrough;
  wire       [7:0]    mac_31_5_io_macOut;
  wire       [7:0]    mac_31_6_io_passthrough;
  wire       [7:0]    mac_31_6_io_macOut;
  wire       [7:0]    mac_31_7_io_passthrough;
  wire       [7:0]    mac_31_7_io_macOut;
  wire       [7:0]    mac_31_8_io_passthrough;
  wire       [7:0]    mac_31_8_io_macOut;
  wire       [7:0]    mac_31_9_io_passthrough;
  wire       [7:0]    mac_31_9_io_macOut;
  wire       [7:0]    mac_31_10_io_passthrough;
  wire       [7:0]    mac_31_10_io_macOut;
  wire       [7:0]    mac_31_11_io_passthrough;
  wire       [7:0]    mac_31_11_io_macOut;
  wire       [7:0]    mac_31_12_io_passthrough;
  wire       [7:0]    mac_31_12_io_macOut;
  wire       [7:0]    mac_31_13_io_passthrough;
  wire       [7:0]    mac_31_13_io_macOut;
  wire       [7:0]    mac_31_14_io_passthrough;
  wire       [7:0]    mac_31_14_io_macOut;
  wire       [7:0]    mac_31_15_io_passthrough;
  wire       [7:0]    mac_31_15_io_macOut;
  wire       [7:0]    mac_31_16_io_passthrough;
  wire       [7:0]    mac_31_16_io_macOut;
  wire       [7:0]    mac_31_17_io_passthrough;
  wire       [7:0]    mac_31_17_io_macOut;
  wire       [7:0]    mac_31_18_io_passthrough;
  wire       [7:0]    mac_31_18_io_macOut;
  wire       [7:0]    mac_31_19_io_passthrough;
  wire       [7:0]    mac_31_19_io_macOut;
  wire       [7:0]    mac_31_20_io_passthrough;
  wire       [7:0]    mac_31_20_io_macOut;
  wire       [7:0]    mac_31_21_io_passthrough;
  wire       [7:0]    mac_31_21_io_macOut;
  wire       [7:0]    mac_31_22_io_passthrough;
  wire       [7:0]    mac_31_22_io_macOut;
  wire       [7:0]    mac_31_23_io_passthrough;
  wire       [7:0]    mac_31_23_io_macOut;
  wire       [7:0]    mac_31_24_io_passthrough;
  wire       [7:0]    mac_31_24_io_macOut;
  wire       [7:0]    mac_31_25_io_passthrough;
  wire       [7:0]    mac_31_25_io_macOut;
  wire       [7:0]    mac_31_26_io_passthrough;
  wire       [7:0]    mac_31_26_io_macOut;
  wire       [7:0]    mac_31_27_io_passthrough;
  wire       [7:0]    mac_31_27_io_macOut;
  wire       [7:0]    mac_31_28_io_passthrough;
  wire       [7:0]    mac_31_28_io_macOut;
  wire       [7:0]    mac_31_29_io_passthrough;
  wire       [7:0]    mac_31_29_io_macOut;
  wire       [7:0]    mac_31_30_io_passthrough;
  wire       [7:0]    mac_31_30_io_macOut;
  wire       [7:0]    mac_31_31_io_passthrough;
  wire       [7:0]    mac_31_31_io_macOut;
  reg        [7:0]    bias_0;
  reg        [7:0]    bias_1;
  reg        [7:0]    bias_2;
  reg        [7:0]    bias_3;
  reg        [7:0]    bias_4;
  reg        [7:0]    bias_5;
  reg        [7:0]    bias_6;
  reg        [7:0]    bias_7;
  reg        [7:0]    bias_8;
  reg        [7:0]    bias_9;
  reg        [7:0]    bias_10;
  reg        [7:0]    bias_11;
  reg        [7:0]    bias_12;
  reg        [7:0]    bias_13;
  reg        [7:0]    bias_14;
  reg        [7:0]    bias_15;
  reg        [7:0]    bias_16;
  reg        [7:0]    bias_17;
  reg        [7:0]    bias_18;
  reg        [7:0]    bias_19;
  reg        [7:0]    bias_20;
  reg        [7:0]    bias_21;
  reg        [7:0]    bias_22;
  reg        [7:0]    bias_23;
  reg        [7:0]    bias_24;
  reg        [7:0]    bias_25;
  reg        [7:0]    bias_26;
  reg        [7:0]    bias_27;
  reg        [7:0]    bias_28;
  reg        [7:0]    bias_29;
  reg        [7:0]    bias_30;
  reg        [7:0]    bias_31;
  reg        [7:0]    io_weight_1_delay_1;
  reg        [7:0]    io_weight_2_delay_1;
  reg        [7:0]    io_weight_2_delay_2;
  reg        [7:0]    io_weight_3_delay_1;
  reg        [7:0]    io_weight_3_delay_2;
  reg        [7:0]    io_weight_3_delay_3;
  reg        [7:0]    io_weight_4_delay_1;
  reg        [7:0]    io_weight_4_delay_2;
  reg        [7:0]    io_weight_4_delay_3;
  reg        [7:0]    io_weight_4_delay_4;
  reg        [7:0]    io_weight_5_delay_1;
  reg        [7:0]    io_weight_5_delay_2;
  reg        [7:0]    io_weight_5_delay_3;
  reg        [7:0]    io_weight_5_delay_4;
  reg        [7:0]    io_weight_5_delay_5;
  reg        [7:0]    io_weight_6_delay_1;
  reg        [7:0]    io_weight_6_delay_2;
  reg        [7:0]    io_weight_6_delay_3;
  reg        [7:0]    io_weight_6_delay_4;
  reg        [7:0]    io_weight_6_delay_5;
  reg        [7:0]    io_weight_6_delay_6;
  reg        [7:0]    io_weight_7_delay_1;
  reg        [7:0]    io_weight_7_delay_2;
  reg        [7:0]    io_weight_7_delay_3;
  reg        [7:0]    io_weight_7_delay_4;
  reg        [7:0]    io_weight_7_delay_5;
  reg        [7:0]    io_weight_7_delay_6;
  reg        [7:0]    io_weight_7_delay_7;
  reg        [7:0]    io_weight_8_delay_1;
  reg        [7:0]    io_weight_8_delay_2;
  reg        [7:0]    io_weight_8_delay_3;
  reg        [7:0]    io_weight_8_delay_4;
  reg        [7:0]    io_weight_8_delay_5;
  reg        [7:0]    io_weight_8_delay_6;
  reg        [7:0]    io_weight_8_delay_7;
  reg        [7:0]    io_weight_8_delay_8;
  reg        [7:0]    io_weight_9_delay_1;
  reg        [7:0]    io_weight_9_delay_2;
  reg        [7:0]    io_weight_9_delay_3;
  reg        [7:0]    io_weight_9_delay_4;
  reg        [7:0]    io_weight_9_delay_5;
  reg        [7:0]    io_weight_9_delay_6;
  reg        [7:0]    io_weight_9_delay_7;
  reg        [7:0]    io_weight_9_delay_8;
  reg        [7:0]    io_weight_9_delay_9;
  reg        [7:0]    io_weight_10_delay_1;
  reg        [7:0]    io_weight_10_delay_2;
  reg        [7:0]    io_weight_10_delay_3;
  reg        [7:0]    io_weight_10_delay_4;
  reg        [7:0]    io_weight_10_delay_5;
  reg        [7:0]    io_weight_10_delay_6;
  reg        [7:0]    io_weight_10_delay_7;
  reg        [7:0]    io_weight_10_delay_8;
  reg        [7:0]    io_weight_10_delay_9;
  reg        [7:0]    io_weight_10_delay_10;
  reg        [7:0]    io_weight_11_delay_1;
  reg        [7:0]    io_weight_11_delay_2;
  reg        [7:0]    io_weight_11_delay_3;
  reg        [7:0]    io_weight_11_delay_4;
  reg        [7:0]    io_weight_11_delay_5;
  reg        [7:0]    io_weight_11_delay_6;
  reg        [7:0]    io_weight_11_delay_7;
  reg        [7:0]    io_weight_11_delay_8;
  reg        [7:0]    io_weight_11_delay_9;
  reg        [7:0]    io_weight_11_delay_10;
  reg        [7:0]    io_weight_11_delay_11;
  reg        [7:0]    io_weight_12_delay_1;
  reg        [7:0]    io_weight_12_delay_2;
  reg        [7:0]    io_weight_12_delay_3;
  reg        [7:0]    io_weight_12_delay_4;
  reg        [7:0]    io_weight_12_delay_5;
  reg        [7:0]    io_weight_12_delay_6;
  reg        [7:0]    io_weight_12_delay_7;
  reg        [7:0]    io_weight_12_delay_8;
  reg        [7:0]    io_weight_12_delay_9;
  reg        [7:0]    io_weight_12_delay_10;
  reg        [7:0]    io_weight_12_delay_11;
  reg        [7:0]    io_weight_12_delay_12;
  reg        [7:0]    io_weight_13_delay_1;
  reg        [7:0]    io_weight_13_delay_2;
  reg        [7:0]    io_weight_13_delay_3;
  reg        [7:0]    io_weight_13_delay_4;
  reg        [7:0]    io_weight_13_delay_5;
  reg        [7:0]    io_weight_13_delay_6;
  reg        [7:0]    io_weight_13_delay_7;
  reg        [7:0]    io_weight_13_delay_8;
  reg        [7:0]    io_weight_13_delay_9;
  reg        [7:0]    io_weight_13_delay_10;
  reg        [7:0]    io_weight_13_delay_11;
  reg        [7:0]    io_weight_13_delay_12;
  reg        [7:0]    io_weight_13_delay_13;
  reg        [7:0]    io_weight_14_delay_1;
  reg        [7:0]    io_weight_14_delay_2;
  reg        [7:0]    io_weight_14_delay_3;
  reg        [7:0]    io_weight_14_delay_4;
  reg        [7:0]    io_weight_14_delay_5;
  reg        [7:0]    io_weight_14_delay_6;
  reg        [7:0]    io_weight_14_delay_7;
  reg        [7:0]    io_weight_14_delay_8;
  reg        [7:0]    io_weight_14_delay_9;
  reg        [7:0]    io_weight_14_delay_10;
  reg        [7:0]    io_weight_14_delay_11;
  reg        [7:0]    io_weight_14_delay_12;
  reg        [7:0]    io_weight_14_delay_13;
  reg        [7:0]    io_weight_14_delay_14;
  reg        [7:0]    io_weight_15_delay_1;
  reg        [7:0]    io_weight_15_delay_2;
  reg        [7:0]    io_weight_15_delay_3;
  reg        [7:0]    io_weight_15_delay_4;
  reg        [7:0]    io_weight_15_delay_5;
  reg        [7:0]    io_weight_15_delay_6;
  reg        [7:0]    io_weight_15_delay_7;
  reg        [7:0]    io_weight_15_delay_8;
  reg        [7:0]    io_weight_15_delay_9;
  reg        [7:0]    io_weight_15_delay_10;
  reg        [7:0]    io_weight_15_delay_11;
  reg        [7:0]    io_weight_15_delay_12;
  reg        [7:0]    io_weight_15_delay_13;
  reg        [7:0]    io_weight_15_delay_14;
  reg        [7:0]    io_weight_15_delay_15;
  reg        [7:0]    io_weight_16_delay_1;
  reg        [7:0]    io_weight_16_delay_2;
  reg        [7:0]    io_weight_16_delay_3;
  reg        [7:0]    io_weight_16_delay_4;
  reg        [7:0]    io_weight_16_delay_5;
  reg        [7:0]    io_weight_16_delay_6;
  reg        [7:0]    io_weight_16_delay_7;
  reg        [7:0]    io_weight_16_delay_8;
  reg        [7:0]    io_weight_16_delay_9;
  reg        [7:0]    io_weight_16_delay_10;
  reg        [7:0]    io_weight_16_delay_11;
  reg        [7:0]    io_weight_16_delay_12;
  reg        [7:0]    io_weight_16_delay_13;
  reg        [7:0]    io_weight_16_delay_14;
  reg        [7:0]    io_weight_16_delay_15;
  reg        [7:0]    io_weight_16_delay_16;
  reg        [7:0]    io_weight_17_delay_1;
  reg        [7:0]    io_weight_17_delay_2;
  reg        [7:0]    io_weight_17_delay_3;
  reg        [7:0]    io_weight_17_delay_4;
  reg        [7:0]    io_weight_17_delay_5;
  reg        [7:0]    io_weight_17_delay_6;
  reg        [7:0]    io_weight_17_delay_7;
  reg        [7:0]    io_weight_17_delay_8;
  reg        [7:0]    io_weight_17_delay_9;
  reg        [7:0]    io_weight_17_delay_10;
  reg        [7:0]    io_weight_17_delay_11;
  reg        [7:0]    io_weight_17_delay_12;
  reg        [7:0]    io_weight_17_delay_13;
  reg        [7:0]    io_weight_17_delay_14;
  reg        [7:0]    io_weight_17_delay_15;
  reg        [7:0]    io_weight_17_delay_16;
  reg        [7:0]    io_weight_17_delay_17;
  reg        [7:0]    io_weight_18_delay_1;
  reg        [7:0]    io_weight_18_delay_2;
  reg        [7:0]    io_weight_18_delay_3;
  reg        [7:0]    io_weight_18_delay_4;
  reg        [7:0]    io_weight_18_delay_5;
  reg        [7:0]    io_weight_18_delay_6;
  reg        [7:0]    io_weight_18_delay_7;
  reg        [7:0]    io_weight_18_delay_8;
  reg        [7:0]    io_weight_18_delay_9;
  reg        [7:0]    io_weight_18_delay_10;
  reg        [7:0]    io_weight_18_delay_11;
  reg        [7:0]    io_weight_18_delay_12;
  reg        [7:0]    io_weight_18_delay_13;
  reg        [7:0]    io_weight_18_delay_14;
  reg        [7:0]    io_weight_18_delay_15;
  reg        [7:0]    io_weight_18_delay_16;
  reg        [7:0]    io_weight_18_delay_17;
  reg        [7:0]    io_weight_18_delay_18;
  reg        [7:0]    io_weight_19_delay_1;
  reg        [7:0]    io_weight_19_delay_2;
  reg        [7:0]    io_weight_19_delay_3;
  reg        [7:0]    io_weight_19_delay_4;
  reg        [7:0]    io_weight_19_delay_5;
  reg        [7:0]    io_weight_19_delay_6;
  reg        [7:0]    io_weight_19_delay_7;
  reg        [7:0]    io_weight_19_delay_8;
  reg        [7:0]    io_weight_19_delay_9;
  reg        [7:0]    io_weight_19_delay_10;
  reg        [7:0]    io_weight_19_delay_11;
  reg        [7:0]    io_weight_19_delay_12;
  reg        [7:0]    io_weight_19_delay_13;
  reg        [7:0]    io_weight_19_delay_14;
  reg        [7:0]    io_weight_19_delay_15;
  reg        [7:0]    io_weight_19_delay_16;
  reg        [7:0]    io_weight_19_delay_17;
  reg        [7:0]    io_weight_19_delay_18;
  reg        [7:0]    io_weight_19_delay_19;
  reg        [7:0]    io_weight_20_delay_1;
  reg        [7:0]    io_weight_20_delay_2;
  reg        [7:0]    io_weight_20_delay_3;
  reg        [7:0]    io_weight_20_delay_4;
  reg        [7:0]    io_weight_20_delay_5;
  reg        [7:0]    io_weight_20_delay_6;
  reg        [7:0]    io_weight_20_delay_7;
  reg        [7:0]    io_weight_20_delay_8;
  reg        [7:0]    io_weight_20_delay_9;
  reg        [7:0]    io_weight_20_delay_10;
  reg        [7:0]    io_weight_20_delay_11;
  reg        [7:0]    io_weight_20_delay_12;
  reg        [7:0]    io_weight_20_delay_13;
  reg        [7:0]    io_weight_20_delay_14;
  reg        [7:0]    io_weight_20_delay_15;
  reg        [7:0]    io_weight_20_delay_16;
  reg        [7:0]    io_weight_20_delay_17;
  reg        [7:0]    io_weight_20_delay_18;
  reg        [7:0]    io_weight_20_delay_19;
  reg        [7:0]    io_weight_20_delay_20;
  reg        [7:0]    io_weight_21_delay_1;
  reg        [7:0]    io_weight_21_delay_2;
  reg        [7:0]    io_weight_21_delay_3;
  reg        [7:0]    io_weight_21_delay_4;
  reg        [7:0]    io_weight_21_delay_5;
  reg        [7:0]    io_weight_21_delay_6;
  reg        [7:0]    io_weight_21_delay_7;
  reg        [7:0]    io_weight_21_delay_8;
  reg        [7:0]    io_weight_21_delay_9;
  reg        [7:0]    io_weight_21_delay_10;
  reg        [7:0]    io_weight_21_delay_11;
  reg        [7:0]    io_weight_21_delay_12;
  reg        [7:0]    io_weight_21_delay_13;
  reg        [7:0]    io_weight_21_delay_14;
  reg        [7:0]    io_weight_21_delay_15;
  reg        [7:0]    io_weight_21_delay_16;
  reg        [7:0]    io_weight_21_delay_17;
  reg        [7:0]    io_weight_21_delay_18;
  reg        [7:0]    io_weight_21_delay_19;
  reg        [7:0]    io_weight_21_delay_20;
  reg        [7:0]    io_weight_21_delay_21;
  reg        [7:0]    io_weight_22_delay_1;
  reg        [7:0]    io_weight_22_delay_2;
  reg        [7:0]    io_weight_22_delay_3;
  reg        [7:0]    io_weight_22_delay_4;
  reg        [7:0]    io_weight_22_delay_5;
  reg        [7:0]    io_weight_22_delay_6;
  reg        [7:0]    io_weight_22_delay_7;
  reg        [7:0]    io_weight_22_delay_8;
  reg        [7:0]    io_weight_22_delay_9;
  reg        [7:0]    io_weight_22_delay_10;
  reg        [7:0]    io_weight_22_delay_11;
  reg        [7:0]    io_weight_22_delay_12;
  reg        [7:0]    io_weight_22_delay_13;
  reg        [7:0]    io_weight_22_delay_14;
  reg        [7:0]    io_weight_22_delay_15;
  reg        [7:0]    io_weight_22_delay_16;
  reg        [7:0]    io_weight_22_delay_17;
  reg        [7:0]    io_weight_22_delay_18;
  reg        [7:0]    io_weight_22_delay_19;
  reg        [7:0]    io_weight_22_delay_20;
  reg        [7:0]    io_weight_22_delay_21;
  reg        [7:0]    io_weight_22_delay_22;
  reg        [7:0]    io_weight_23_delay_1;
  reg        [7:0]    io_weight_23_delay_2;
  reg        [7:0]    io_weight_23_delay_3;
  reg        [7:0]    io_weight_23_delay_4;
  reg        [7:0]    io_weight_23_delay_5;
  reg        [7:0]    io_weight_23_delay_6;
  reg        [7:0]    io_weight_23_delay_7;
  reg        [7:0]    io_weight_23_delay_8;
  reg        [7:0]    io_weight_23_delay_9;
  reg        [7:0]    io_weight_23_delay_10;
  reg        [7:0]    io_weight_23_delay_11;
  reg        [7:0]    io_weight_23_delay_12;
  reg        [7:0]    io_weight_23_delay_13;
  reg        [7:0]    io_weight_23_delay_14;
  reg        [7:0]    io_weight_23_delay_15;
  reg        [7:0]    io_weight_23_delay_16;
  reg        [7:0]    io_weight_23_delay_17;
  reg        [7:0]    io_weight_23_delay_18;
  reg        [7:0]    io_weight_23_delay_19;
  reg        [7:0]    io_weight_23_delay_20;
  reg        [7:0]    io_weight_23_delay_21;
  reg        [7:0]    io_weight_23_delay_22;
  reg        [7:0]    io_weight_23_delay_23;
  reg        [7:0]    io_weight_24_delay_1;
  reg        [7:0]    io_weight_24_delay_2;
  reg        [7:0]    io_weight_24_delay_3;
  reg        [7:0]    io_weight_24_delay_4;
  reg        [7:0]    io_weight_24_delay_5;
  reg        [7:0]    io_weight_24_delay_6;
  reg        [7:0]    io_weight_24_delay_7;
  reg        [7:0]    io_weight_24_delay_8;
  reg        [7:0]    io_weight_24_delay_9;
  reg        [7:0]    io_weight_24_delay_10;
  reg        [7:0]    io_weight_24_delay_11;
  reg        [7:0]    io_weight_24_delay_12;
  reg        [7:0]    io_weight_24_delay_13;
  reg        [7:0]    io_weight_24_delay_14;
  reg        [7:0]    io_weight_24_delay_15;
  reg        [7:0]    io_weight_24_delay_16;
  reg        [7:0]    io_weight_24_delay_17;
  reg        [7:0]    io_weight_24_delay_18;
  reg        [7:0]    io_weight_24_delay_19;
  reg        [7:0]    io_weight_24_delay_20;
  reg        [7:0]    io_weight_24_delay_21;
  reg        [7:0]    io_weight_24_delay_22;
  reg        [7:0]    io_weight_24_delay_23;
  reg        [7:0]    io_weight_24_delay_24;
  reg        [7:0]    io_weight_25_delay_1;
  reg        [7:0]    io_weight_25_delay_2;
  reg        [7:0]    io_weight_25_delay_3;
  reg        [7:0]    io_weight_25_delay_4;
  reg        [7:0]    io_weight_25_delay_5;
  reg        [7:0]    io_weight_25_delay_6;
  reg        [7:0]    io_weight_25_delay_7;
  reg        [7:0]    io_weight_25_delay_8;
  reg        [7:0]    io_weight_25_delay_9;
  reg        [7:0]    io_weight_25_delay_10;
  reg        [7:0]    io_weight_25_delay_11;
  reg        [7:0]    io_weight_25_delay_12;
  reg        [7:0]    io_weight_25_delay_13;
  reg        [7:0]    io_weight_25_delay_14;
  reg        [7:0]    io_weight_25_delay_15;
  reg        [7:0]    io_weight_25_delay_16;
  reg        [7:0]    io_weight_25_delay_17;
  reg        [7:0]    io_weight_25_delay_18;
  reg        [7:0]    io_weight_25_delay_19;
  reg        [7:0]    io_weight_25_delay_20;
  reg        [7:0]    io_weight_25_delay_21;
  reg        [7:0]    io_weight_25_delay_22;
  reg        [7:0]    io_weight_25_delay_23;
  reg        [7:0]    io_weight_25_delay_24;
  reg        [7:0]    io_weight_25_delay_25;
  reg        [7:0]    io_weight_26_delay_1;
  reg        [7:0]    io_weight_26_delay_2;
  reg        [7:0]    io_weight_26_delay_3;
  reg        [7:0]    io_weight_26_delay_4;
  reg        [7:0]    io_weight_26_delay_5;
  reg        [7:0]    io_weight_26_delay_6;
  reg        [7:0]    io_weight_26_delay_7;
  reg        [7:0]    io_weight_26_delay_8;
  reg        [7:0]    io_weight_26_delay_9;
  reg        [7:0]    io_weight_26_delay_10;
  reg        [7:0]    io_weight_26_delay_11;
  reg        [7:0]    io_weight_26_delay_12;
  reg        [7:0]    io_weight_26_delay_13;
  reg        [7:0]    io_weight_26_delay_14;
  reg        [7:0]    io_weight_26_delay_15;
  reg        [7:0]    io_weight_26_delay_16;
  reg        [7:0]    io_weight_26_delay_17;
  reg        [7:0]    io_weight_26_delay_18;
  reg        [7:0]    io_weight_26_delay_19;
  reg        [7:0]    io_weight_26_delay_20;
  reg        [7:0]    io_weight_26_delay_21;
  reg        [7:0]    io_weight_26_delay_22;
  reg        [7:0]    io_weight_26_delay_23;
  reg        [7:0]    io_weight_26_delay_24;
  reg        [7:0]    io_weight_26_delay_25;
  reg        [7:0]    io_weight_26_delay_26;
  reg        [7:0]    io_weight_27_delay_1;
  reg        [7:0]    io_weight_27_delay_2;
  reg        [7:0]    io_weight_27_delay_3;
  reg        [7:0]    io_weight_27_delay_4;
  reg        [7:0]    io_weight_27_delay_5;
  reg        [7:0]    io_weight_27_delay_6;
  reg        [7:0]    io_weight_27_delay_7;
  reg        [7:0]    io_weight_27_delay_8;
  reg        [7:0]    io_weight_27_delay_9;
  reg        [7:0]    io_weight_27_delay_10;
  reg        [7:0]    io_weight_27_delay_11;
  reg        [7:0]    io_weight_27_delay_12;
  reg        [7:0]    io_weight_27_delay_13;
  reg        [7:0]    io_weight_27_delay_14;
  reg        [7:0]    io_weight_27_delay_15;
  reg        [7:0]    io_weight_27_delay_16;
  reg        [7:0]    io_weight_27_delay_17;
  reg        [7:0]    io_weight_27_delay_18;
  reg        [7:0]    io_weight_27_delay_19;
  reg        [7:0]    io_weight_27_delay_20;
  reg        [7:0]    io_weight_27_delay_21;
  reg        [7:0]    io_weight_27_delay_22;
  reg        [7:0]    io_weight_27_delay_23;
  reg        [7:0]    io_weight_27_delay_24;
  reg        [7:0]    io_weight_27_delay_25;
  reg        [7:0]    io_weight_27_delay_26;
  reg        [7:0]    io_weight_27_delay_27;
  reg        [7:0]    io_weight_28_delay_1;
  reg        [7:0]    io_weight_28_delay_2;
  reg        [7:0]    io_weight_28_delay_3;
  reg        [7:0]    io_weight_28_delay_4;
  reg        [7:0]    io_weight_28_delay_5;
  reg        [7:0]    io_weight_28_delay_6;
  reg        [7:0]    io_weight_28_delay_7;
  reg        [7:0]    io_weight_28_delay_8;
  reg        [7:0]    io_weight_28_delay_9;
  reg        [7:0]    io_weight_28_delay_10;
  reg        [7:0]    io_weight_28_delay_11;
  reg        [7:0]    io_weight_28_delay_12;
  reg        [7:0]    io_weight_28_delay_13;
  reg        [7:0]    io_weight_28_delay_14;
  reg        [7:0]    io_weight_28_delay_15;
  reg        [7:0]    io_weight_28_delay_16;
  reg        [7:0]    io_weight_28_delay_17;
  reg        [7:0]    io_weight_28_delay_18;
  reg        [7:0]    io_weight_28_delay_19;
  reg        [7:0]    io_weight_28_delay_20;
  reg        [7:0]    io_weight_28_delay_21;
  reg        [7:0]    io_weight_28_delay_22;
  reg        [7:0]    io_weight_28_delay_23;
  reg        [7:0]    io_weight_28_delay_24;
  reg        [7:0]    io_weight_28_delay_25;
  reg        [7:0]    io_weight_28_delay_26;
  reg        [7:0]    io_weight_28_delay_27;
  reg        [7:0]    io_weight_28_delay_28;
  reg        [7:0]    io_weight_29_delay_1;
  reg        [7:0]    io_weight_29_delay_2;
  reg        [7:0]    io_weight_29_delay_3;
  reg        [7:0]    io_weight_29_delay_4;
  reg        [7:0]    io_weight_29_delay_5;
  reg        [7:0]    io_weight_29_delay_6;
  reg        [7:0]    io_weight_29_delay_7;
  reg        [7:0]    io_weight_29_delay_8;
  reg        [7:0]    io_weight_29_delay_9;
  reg        [7:0]    io_weight_29_delay_10;
  reg        [7:0]    io_weight_29_delay_11;
  reg        [7:0]    io_weight_29_delay_12;
  reg        [7:0]    io_weight_29_delay_13;
  reg        [7:0]    io_weight_29_delay_14;
  reg        [7:0]    io_weight_29_delay_15;
  reg        [7:0]    io_weight_29_delay_16;
  reg        [7:0]    io_weight_29_delay_17;
  reg        [7:0]    io_weight_29_delay_18;
  reg        [7:0]    io_weight_29_delay_19;
  reg        [7:0]    io_weight_29_delay_20;
  reg        [7:0]    io_weight_29_delay_21;
  reg        [7:0]    io_weight_29_delay_22;
  reg        [7:0]    io_weight_29_delay_23;
  reg        [7:0]    io_weight_29_delay_24;
  reg        [7:0]    io_weight_29_delay_25;
  reg        [7:0]    io_weight_29_delay_26;
  reg        [7:0]    io_weight_29_delay_27;
  reg        [7:0]    io_weight_29_delay_28;
  reg        [7:0]    io_weight_29_delay_29;
  reg        [7:0]    io_weight_30_delay_1;
  reg        [7:0]    io_weight_30_delay_2;
  reg        [7:0]    io_weight_30_delay_3;
  reg        [7:0]    io_weight_30_delay_4;
  reg        [7:0]    io_weight_30_delay_5;
  reg        [7:0]    io_weight_30_delay_6;
  reg        [7:0]    io_weight_30_delay_7;
  reg        [7:0]    io_weight_30_delay_8;
  reg        [7:0]    io_weight_30_delay_9;
  reg        [7:0]    io_weight_30_delay_10;
  reg        [7:0]    io_weight_30_delay_11;
  reg        [7:0]    io_weight_30_delay_12;
  reg        [7:0]    io_weight_30_delay_13;
  reg        [7:0]    io_weight_30_delay_14;
  reg        [7:0]    io_weight_30_delay_15;
  reg        [7:0]    io_weight_30_delay_16;
  reg        [7:0]    io_weight_30_delay_17;
  reg        [7:0]    io_weight_30_delay_18;
  reg        [7:0]    io_weight_30_delay_19;
  reg        [7:0]    io_weight_30_delay_20;
  reg        [7:0]    io_weight_30_delay_21;
  reg        [7:0]    io_weight_30_delay_22;
  reg        [7:0]    io_weight_30_delay_23;
  reg        [7:0]    io_weight_30_delay_24;
  reg        [7:0]    io_weight_30_delay_25;
  reg        [7:0]    io_weight_30_delay_26;
  reg        [7:0]    io_weight_30_delay_27;
  reg        [7:0]    io_weight_30_delay_28;
  reg        [7:0]    io_weight_30_delay_29;
  reg        [7:0]    io_weight_30_delay_30;
  reg        [7:0]    io_weight_31_delay_1;
  reg        [7:0]    io_weight_31_delay_2;
  reg        [7:0]    io_weight_31_delay_3;
  reg        [7:0]    io_weight_31_delay_4;
  reg        [7:0]    io_weight_31_delay_5;
  reg        [7:0]    io_weight_31_delay_6;
  reg        [7:0]    io_weight_31_delay_7;
  reg        [7:0]    io_weight_31_delay_8;
  reg        [7:0]    io_weight_31_delay_9;
  reg        [7:0]    io_weight_31_delay_10;
  reg        [7:0]    io_weight_31_delay_11;
  reg        [7:0]    io_weight_31_delay_12;
  reg        [7:0]    io_weight_31_delay_13;
  reg        [7:0]    io_weight_31_delay_14;
  reg        [7:0]    io_weight_31_delay_15;
  reg        [7:0]    io_weight_31_delay_16;
  reg        [7:0]    io_weight_31_delay_17;
  reg        [7:0]    io_weight_31_delay_18;
  reg        [7:0]    io_weight_31_delay_19;
  reg        [7:0]    io_weight_31_delay_20;
  reg        [7:0]    io_weight_31_delay_21;
  reg        [7:0]    io_weight_31_delay_22;
  reg        [7:0]    io_weight_31_delay_23;
  reg        [7:0]    io_weight_31_delay_24;
  reg        [7:0]    io_weight_31_delay_25;
  reg        [7:0]    io_weight_31_delay_26;
  reg        [7:0]    io_weight_31_delay_27;
  reg        [7:0]    io_weight_31_delay_28;
  reg        [7:0]    io_weight_31_delay_29;
  reg        [7:0]    io_weight_31_delay_30;
  reg        [7:0]    io_weight_31_delay_31;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_9;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_10;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_11;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_12;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_13;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_14;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_15;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_16;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_17;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_18;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_19;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_20;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_21;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_22;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_23;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_24;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_25;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_26;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_27;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_28;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_29;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_30;
  reg        [7:0]    toplevel_mac_0_31_io_macOut_delay_31;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_9;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_10;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_11;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_12;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_13;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_14;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_15;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_16;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_17;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_18;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_19;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_20;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_21;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_22;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_23;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_24;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_25;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_26;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_27;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_28;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_29;
  reg        [7:0]    toplevel_mac_1_31_io_macOut_delay_30;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_9;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_10;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_11;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_12;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_13;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_14;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_15;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_16;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_17;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_18;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_19;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_20;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_21;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_22;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_23;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_24;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_25;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_26;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_27;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_28;
  reg        [7:0]    toplevel_mac_2_31_io_macOut_delay_29;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_9;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_10;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_11;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_12;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_13;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_14;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_15;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_16;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_17;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_18;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_19;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_20;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_21;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_22;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_23;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_24;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_25;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_26;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_27;
  reg        [7:0]    toplevel_mac_3_31_io_macOut_delay_28;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_9;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_10;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_11;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_12;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_13;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_14;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_15;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_16;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_17;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_18;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_19;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_20;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_21;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_22;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_23;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_24;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_25;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_26;
  reg        [7:0]    toplevel_mac_4_31_io_macOut_delay_27;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_9;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_10;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_11;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_12;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_13;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_14;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_15;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_16;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_17;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_18;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_19;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_20;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_21;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_22;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_23;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_24;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_25;
  reg        [7:0]    toplevel_mac_5_31_io_macOut_delay_26;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_9;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_10;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_11;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_12;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_13;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_14;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_15;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_16;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_17;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_18;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_19;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_20;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_21;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_22;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_23;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_24;
  reg        [7:0]    toplevel_mac_6_31_io_macOut_delay_25;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_9;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_10;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_11;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_12;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_13;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_14;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_15;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_16;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_17;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_18;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_19;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_20;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_21;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_22;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_23;
  reg        [7:0]    toplevel_mac_7_31_io_macOut_delay_24;
  reg        [7:0]    toplevel_mac_8_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_8_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_8_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_8_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_8_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_8_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_8_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_8_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_8_31_io_macOut_delay_9;
  reg        [7:0]    toplevel_mac_8_31_io_macOut_delay_10;
  reg        [7:0]    toplevel_mac_8_31_io_macOut_delay_11;
  reg        [7:0]    toplevel_mac_8_31_io_macOut_delay_12;
  reg        [7:0]    toplevel_mac_8_31_io_macOut_delay_13;
  reg        [7:0]    toplevel_mac_8_31_io_macOut_delay_14;
  reg        [7:0]    toplevel_mac_8_31_io_macOut_delay_15;
  reg        [7:0]    toplevel_mac_8_31_io_macOut_delay_16;
  reg        [7:0]    toplevel_mac_8_31_io_macOut_delay_17;
  reg        [7:0]    toplevel_mac_8_31_io_macOut_delay_18;
  reg        [7:0]    toplevel_mac_8_31_io_macOut_delay_19;
  reg        [7:0]    toplevel_mac_8_31_io_macOut_delay_20;
  reg        [7:0]    toplevel_mac_8_31_io_macOut_delay_21;
  reg        [7:0]    toplevel_mac_8_31_io_macOut_delay_22;
  reg        [7:0]    toplevel_mac_8_31_io_macOut_delay_23;
  reg        [7:0]    toplevel_mac_9_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_9_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_9_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_9_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_9_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_9_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_9_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_9_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_9_31_io_macOut_delay_9;
  reg        [7:0]    toplevel_mac_9_31_io_macOut_delay_10;
  reg        [7:0]    toplevel_mac_9_31_io_macOut_delay_11;
  reg        [7:0]    toplevel_mac_9_31_io_macOut_delay_12;
  reg        [7:0]    toplevel_mac_9_31_io_macOut_delay_13;
  reg        [7:0]    toplevel_mac_9_31_io_macOut_delay_14;
  reg        [7:0]    toplevel_mac_9_31_io_macOut_delay_15;
  reg        [7:0]    toplevel_mac_9_31_io_macOut_delay_16;
  reg        [7:0]    toplevel_mac_9_31_io_macOut_delay_17;
  reg        [7:0]    toplevel_mac_9_31_io_macOut_delay_18;
  reg        [7:0]    toplevel_mac_9_31_io_macOut_delay_19;
  reg        [7:0]    toplevel_mac_9_31_io_macOut_delay_20;
  reg        [7:0]    toplevel_mac_9_31_io_macOut_delay_21;
  reg        [7:0]    toplevel_mac_9_31_io_macOut_delay_22;
  reg        [7:0]    toplevel_mac_10_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_10_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_10_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_10_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_10_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_10_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_10_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_10_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_10_31_io_macOut_delay_9;
  reg        [7:0]    toplevel_mac_10_31_io_macOut_delay_10;
  reg        [7:0]    toplevel_mac_10_31_io_macOut_delay_11;
  reg        [7:0]    toplevel_mac_10_31_io_macOut_delay_12;
  reg        [7:0]    toplevel_mac_10_31_io_macOut_delay_13;
  reg        [7:0]    toplevel_mac_10_31_io_macOut_delay_14;
  reg        [7:0]    toplevel_mac_10_31_io_macOut_delay_15;
  reg        [7:0]    toplevel_mac_10_31_io_macOut_delay_16;
  reg        [7:0]    toplevel_mac_10_31_io_macOut_delay_17;
  reg        [7:0]    toplevel_mac_10_31_io_macOut_delay_18;
  reg        [7:0]    toplevel_mac_10_31_io_macOut_delay_19;
  reg        [7:0]    toplevel_mac_10_31_io_macOut_delay_20;
  reg        [7:0]    toplevel_mac_10_31_io_macOut_delay_21;
  reg        [7:0]    toplevel_mac_11_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_11_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_11_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_11_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_11_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_11_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_11_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_11_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_11_31_io_macOut_delay_9;
  reg        [7:0]    toplevel_mac_11_31_io_macOut_delay_10;
  reg        [7:0]    toplevel_mac_11_31_io_macOut_delay_11;
  reg        [7:0]    toplevel_mac_11_31_io_macOut_delay_12;
  reg        [7:0]    toplevel_mac_11_31_io_macOut_delay_13;
  reg        [7:0]    toplevel_mac_11_31_io_macOut_delay_14;
  reg        [7:0]    toplevel_mac_11_31_io_macOut_delay_15;
  reg        [7:0]    toplevel_mac_11_31_io_macOut_delay_16;
  reg        [7:0]    toplevel_mac_11_31_io_macOut_delay_17;
  reg        [7:0]    toplevel_mac_11_31_io_macOut_delay_18;
  reg        [7:0]    toplevel_mac_11_31_io_macOut_delay_19;
  reg        [7:0]    toplevel_mac_11_31_io_macOut_delay_20;
  reg        [7:0]    toplevel_mac_12_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_12_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_12_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_12_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_12_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_12_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_12_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_12_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_12_31_io_macOut_delay_9;
  reg        [7:0]    toplevel_mac_12_31_io_macOut_delay_10;
  reg        [7:0]    toplevel_mac_12_31_io_macOut_delay_11;
  reg        [7:0]    toplevel_mac_12_31_io_macOut_delay_12;
  reg        [7:0]    toplevel_mac_12_31_io_macOut_delay_13;
  reg        [7:0]    toplevel_mac_12_31_io_macOut_delay_14;
  reg        [7:0]    toplevel_mac_12_31_io_macOut_delay_15;
  reg        [7:0]    toplevel_mac_12_31_io_macOut_delay_16;
  reg        [7:0]    toplevel_mac_12_31_io_macOut_delay_17;
  reg        [7:0]    toplevel_mac_12_31_io_macOut_delay_18;
  reg        [7:0]    toplevel_mac_12_31_io_macOut_delay_19;
  reg        [7:0]    toplevel_mac_13_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_13_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_13_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_13_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_13_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_13_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_13_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_13_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_13_31_io_macOut_delay_9;
  reg        [7:0]    toplevel_mac_13_31_io_macOut_delay_10;
  reg        [7:0]    toplevel_mac_13_31_io_macOut_delay_11;
  reg        [7:0]    toplevel_mac_13_31_io_macOut_delay_12;
  reg        [7:0]    toplevel_mac_13_31_io_macOut_delay_13;
  reg        [7:0]    toplevel_mac_13_31_io_macOut_delay_14;
  reg        [7:0]    toplevel_mac_13_31_io_macOut_delay_15;
  reg        [7:0]    toplevel_mac_13_31_io_macOut_delay_16;
  reg        [7:0]    toplevel_mac_13_31_io_macOut_delay_17;
  reg        [7:0]    toplevel_mac_13_31_io_macOut_delay_18;
  reg        [7:0]    toplevel_mac_14_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_14_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_14_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_14_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_14_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_14_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_14_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_14_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_14_31_io_macOut_delay_9;
  reg        [7:0]    toplevel_mac_14_31_io_macOut_delay_10;
  reg        [7:0]    toplevel_mac_14_31_io_macOut_delay_11;
  reg        [7:0]    toplevel_mac_14_31_io_macOut_delay_12;
  reg        [7:0]    toplevel_mac_14_31_io_macOut_delay_13;
  reg        [7:0]    toplevel_mac_14_31_io_macOut_delay_14;
  reg        [7:0]    toplevel_mac_14_31_io_macOut_delay_15;
  reg        [7:0]    toplevel_mac_14_31_io_macOut_delay_16;
  reg        [7:0]    toplevel_mac_14_31_io_macOut_delay_17;
  reg        [7:0]    toplevel_mac_15_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_15_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_15_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_15_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_15_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_15_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_15_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_15_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_15_31_io_macOut_delay_9;
  reg        [7:0]    toplevel_mac_15_31_io_macOut_delay_10;
  reg        [7:0]    toplevel_mac_15_31_io_macOut_delay_11;
  reg        [7:0]    toplevel_mac_15_31_io_macOut_delay_12;
  reg        [7:0]    toplevel_mac_15_31_io_macOut_delay_13;
  reg        [7:0]    toplevel_mac_15_31_io_macOut_delay_14;
  reg        [7:0]    toplevel_mac_15_31_io_macOut_delay_15;
  reg        [7:0]    toplevel_mac_15_31_io_macOut_delay_16;
  reg        [7:0]    toplevel_mac_16_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_16_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_16_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_16_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_16_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_16_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_16_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_16_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_16_31_io_macOut_delay_9;
  reg        [7:0]    toplevel_mac_16_31_io_macOut_delay_10;
  reg        [7:0]    toplevel_mac_16_31_io_macOut_delay_11;
  reg        [7:0]    toplevel_mac_16_31_io_macOut_delay_12;
  reg        [7:0]    toplevel_mac_16_31_io_macOut_delay_13;
  reg        [7:0]    toplevel_mac_16_31_io_macOut_delay_14;
  reg        [7:0]    toplevel_mac_16_31_io_macOut_delay_15;
  reg        [7:0]    toplevel_mac_17_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_17_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_17_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_17_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_17_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_17_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_17_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_17_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_17_31_io_macOut_delay_9;
  reg        [7:0]    toplevel_mac_17_31_io_macOut_delay_10;
  reg        [7:0]    toplevel_mac_17_31_io_macOut_delay_11;
  reg        [7:0]    toplevel_mac_17_31_io_macOut_delay_12;
  reg        [7:0]    toplevel_mac_17_31_io_macOut_delay_13;
  reg        [7:0]    toplevel_mac_17_31_io_macOut_delay_14;
  reg        [7:0]    toplevel_mac_18_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_18_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_18_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_18_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_18_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_18_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_18_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_18_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_18_31_io_macOut_delay_9;
  reg        [7:0]    toplevel_mac_18_31_io_macOut_delay_10;
  reg        [7:0]    toplevel_mac_18_31_io_macOut_delay_11;
  reg        [7:0]    toplevel_mac_18_31_io_macOut_delay_12;
  reg        [7:0]    toplevel_mac_18_31_io_macOut_delay_13;
  reg        [7:0]    toplevel_mac_19_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_19_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_19_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_19_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_19_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_19_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_19_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_19_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_19_31_io_macOut_delay_9;
  reg        [7:0]    toplevel_mac_19_31_io_macOut_delay_10;
  reg        [7:0]    toplevel_mac_19_31_io_macOut_delay_11;
  reg        [7:0]    toplevel_mac_19_31_io_macOut_delay_12;
  reg        [7:0]    toplevel_mac_20_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_20_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_20_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_20_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_20_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_20_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_20_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_20_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_20_31_io_macOut_delay_9;
  reg        [7:0]    toplevel_mac_20_31_io_macOut_delay_10;
  reg        [7:0]    toplevel_mac_20_31_io_macOut_delay_11;
  reg        [7:0]    toplevel_mac_21_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_21_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_21_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_21_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_21_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_21_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_21_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_21_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_21_31_io_macOut_delay_9;
  reg        [7:0]    toplevel_mac_21_31_io_macOut_delay_10;
  reg        [7:0]    toplevel_mac_22_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_22_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_22_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_22_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_22_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_22_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_22_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_22_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_22_31_io_macOut_delay_9;
  reg        [7:0]    toplevel_mac_23_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_23_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_23_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_23_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_23_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_23_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_23_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_23_31_io_macOut_delay_8;
  reg        [7:0]    toplevel_mac_24_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_24_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_24_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_24_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_24_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_24_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_24_31_io_macOut_delay_7;
  reg        [7:0]    toplevel_mac_25_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_25_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_25_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_25_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_25_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_25_31_io_macOut_delay_6;
  reg        [7:0]    toplevel_mac_26_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_26_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_26_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_26_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_26_31_io_macOut_delay_5;
  reg        [7:0]    toplevel_mac_27_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_27_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_27_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_27_31_io_macOut_delay_4;
  reg        [7:0]    toplevel_mac_28_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_28_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_28_31_io_macOut_delay_3;
  reg        [7:0]    toplevel_mac_29_31_io_macOut_delay_1;
  reg        [7:0]    toplevel_mac_29_31_io_macOut_delay_2;
  reg        [7:0]    toplevel_mac_30_31_io_macOut_delay_1;

  MAC mac_0_0 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (io_weight_0[7:0]           ), //i
    .io_addInput    (bias_0[7:0]                ), //i
    .io_passthrough (mac_0_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_0_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_1 mac_0_1 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (io_weight_1_delay_1[7:0]   ), //i
    .io_addInput    (mac_0_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_1_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_2 mac_0_2 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (io_weight_2_delay_2[7:0]   ), //i
    .io_addInput    (mac_0_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_2_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_3 mac_0_3 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (io_weight_3_delay_3[7:0]   ), //i
    .io_addInput    (mac_0_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_3_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_4 mac_0_4 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (io_weight_4_delay_4[7:0]   ), //i
    .io_addInput    (mac_0_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_4_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_5 mac_0_5 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (io_weight_5_delay_5[7:0]   ), //i
    .io_addInput    (mac_0_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_5_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_6 mac_0_6 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (io_weight_6_delay_6[7:0]   ), //i
    .io_addInput    (mac_0_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_6_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_7 mac_0_7 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (io_weight_7_delay_7[7:0]   ), //i
    .io_addInput    (mac_0_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_7_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_8 mac_0_8 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (io_weight_8_delay_8[7:0]   ), //i
    .io_addInput    (mac_0_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_8_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_9 mac_0_9 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (io_weight_9_delay_9[7:0]   ), //i
    .io_addInput    (mac_0_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_9_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_10 mac_0_10 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (io_weight_10_delay_10[7:0]  ), //i
    .io_addInput    (mac_0_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_0_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_10_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_11 mac_0_11 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (io_weight_11_delay_11[7:0]  ), //i
    .io_addInput    (mac_0_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_11_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_12 mac_0_12 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (io_weight_12_delay_12[7:0]  ), //i
    .io_addInput    (mac_0_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_12_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_13 mac_0_13 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (io_weight_13_delay_13[7:0]  ), //i
    .io_addInput    (mac_0_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_13_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_14 mac_0_14 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (io_weight_14_delay_14[7:0]  ), //i
    .io_addInput    (mac_0_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_14_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_15 mac_0_15 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (io_weight_15_delay_15[7:0]  ), //i
    .io_addInput    (mac_0_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_15_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_16 mac_0_16 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (io_weight_16_delay_16[7:0]  ), //i
    .io_addInput    (mac_0_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_16_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_17 mac_0_17 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (io_weight_17_delay_17[7:0]  ), //i
    .io_addInput    (mac_0_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_17_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_18 mac_0_18 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (io_weight_18_delay_18[7:0]  ), //i
    .io_addInput    (mac_0_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_18_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_19 mac_0_19 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (io_weight_19_delay_19[7:0]  ), //i
    .io_addInput    (mac_0_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_19_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_20 mac_0_20 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (io_weight_20_delay_20[7:0]  ), //i
    .io_addInput    (mac_0_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_20_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_21 mac_0_21 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (io_weight_21_delay_21[7:0]  ), //i
    .io_addInput    (mac_0_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_21_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_22 mac_0_22 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (io_weight_22_delay_22[7:0]  ), //i
    .io_addInput    (mac_0_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_22_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_23 mac_0_23 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (io_weight_23_delay_23[7:0]  ), //i
    .io_addInput    (mac_0_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_23_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_24 mac_0_24 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (io_weight_24_delay_24[7:0]  ), //i
    .io_addInput    (mac_0_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_24_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_25 mac_0_25 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (io_weight_25_delay_25[7:0]  ), //i
    .io_addInput    (mac_0_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_25_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_26 mac_0_26 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (io_weight_26_delay_26[7:0]  ), //i
    .io_addInput    (mac_0_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_26_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_27 mac_0_27 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (io_weight_27_delay_27[7:0]  ), //i
    .io_addInput    (mac_0_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_27_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_28 mac_0_28 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (io_weight_28_delay_28[7:0]  ), //i
    .io_addInput    (mac_0_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_28_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_29 mac_0_29 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (io_weight_29_delay_29[7:0]  ), //i
    .io_addInput    (mac_0_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_29_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_30 mac_0_30 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (io_weight_30_delay_30[7:0]  ), //i
    .io_addInput    (mac_0_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_30_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_31 mac_0_31 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (io_weight_31_delay_31[7:0]  ), //i
    .io_addInput    (mac_0_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_0_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_0_31_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_32 mac_1_0 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_0_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_1[7:0]                ), //i
    .io_passthrough (mac_1_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_0_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_33 mac_1_1 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_0_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_1_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_34 mac_1_2 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_0_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_2_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_35 mac_1_3 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_0_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_3_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_36 mac_1_4 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_0_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_4_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_37 mac_1_5 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_0_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_5_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_38 mac_1_6 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_0_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_6_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_39 mac_1_7 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_0_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_7_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_40 mac_1_8 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_0_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_8_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_41 mac_1_9 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_0_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_9_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_42 mac_1_10 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_0_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_1_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_10_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_43 mac_1_11 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_0_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_11_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_44 mac_1_12 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_0_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_12_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_45 mac_1_13 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_0_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_13_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_46 mac_1_14 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_0_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_14_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_47 mac_1_15 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_0_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_15_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_48 mac_1_16 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_0_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_16_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_49 mac_1_17 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_0_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_17_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_50 mac_1_18 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_0_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_18_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_51 mac_1_19 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_0_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_19_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_52 mac_1_20 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_0_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_20_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_53 mac_1_21 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_0_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_21_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_54 mac_1_22 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_0_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_22_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_55 mac_1_23 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_0_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_23_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_56 mac_1_24 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_0_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_24_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_57 mac_1_25 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_0_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_25_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_58 mac_1_26 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_0_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_26_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_59 mac_1_27 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_0_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_27_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_60 mac_1_28 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_0_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_28_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_61 mac_1_29 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_0_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_29_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_62 mac_1_30 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_0_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_30_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_63 mac_1_31 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_0_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_1_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_1_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_1_31_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_64 mac_2_0 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_1_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_2[7:0]                ), //i
    .io_passthrough (mac_2_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_0_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_65 mac_2_1 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_1_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_1_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_66 mac_2_2 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_1_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_2_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_67 mac_2_3 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_1_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_3_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_68 mac_2_4 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_1_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_4_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_69 mac_2_5 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_1_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_5_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_70 mac_2_6 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_1_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_6_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_71 mac_2_7 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_1_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_7_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_72 mac_2_8 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_1_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_8_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_73 mac_2_9 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_1_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_9_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_74 mac_2_10 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_1_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_2_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_10_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_75 mac_2_11 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_1_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_11_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_76 mac_2_12 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_1_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_12_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_77 mac_2_13 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_1_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_13_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_78 mac_2_14 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_1_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_14_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_79 mac_2_15 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_1_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_15_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_80 mac_2_16 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_1_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_16_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_81 mac_2_17 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_1_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_17_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_82 mac_2_18 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_1_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_18_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_83 mac_2_19 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_1_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_19_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_84 mac_2_20 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_1_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_20_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_85 mac_2_21 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_1_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_21_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_86 mac_2_22 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_1_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_22_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_87 mac_2_23 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_1_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_23_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_88 mac_2_24 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_1_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_24_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_89 mac_2_25 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_1_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_25_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_90 mac_2_26 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_1_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_26_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_91 mac_2_27 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_1_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_27_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_92 mac_2_28 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_1_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_28_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_93 mac_2_29 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_1_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_29_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_94 mac_2_30 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_1_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_30_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_95 mac_2_31 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_1_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_2_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_2_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_2_31_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_96 mac_3_0 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_2_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_3[7:0]                ), //i
    .io_passthrough (mac_3_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_0_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_97 mac_3_1 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_2_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_1_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_98 mac_3_2 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_2_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_2_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_99 mac_3_3 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_2_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_3_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_100 mac_3_4 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_2_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_4_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_101 mac_3_5 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_2_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_5_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_102 mac_3_6 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_2_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_6_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_103 mac_3_7 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_2_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_7_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_104 mac_3_8 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_2_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_8_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_105 mac_3_9 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_2_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_9_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_106 mac_3_10 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_2_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_3_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_10_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_107 mac_3_11 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_2_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_11_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_108 mac_3_12 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_2_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_12_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_109 mac_3_13 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_2_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_13_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_110 mac_3_14 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_2_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_14_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_111 mac_3_15 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_2_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_15_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_112 mac_3_16 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_2_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_16_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_113 mac_3_17 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_2_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_17_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_114 mac_3_18 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_2_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_18_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_115 mac_3_19 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_2_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_19_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_116 mac_3_20 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_2_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_20_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_117 mac_3_21 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_2_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_21_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_118 mac_3_22 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_2_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_22_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_119 mac_3_23 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_2_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_23_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_120 mac_3_24 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_2_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_24_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_121 mac_3_25 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_2_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_25_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_122 mac_3_26 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_2_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_26_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_123 mac_3_27 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_2_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_27_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_124 mac_3_28 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_2_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_28_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_125 mac_3_29 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_2_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_29_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_126 mac_3_30 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_2_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_30_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_127 mac_3_31 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_2_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_3_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_3_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_3_31_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_128 mac_4_0 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_3_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_4[7:0]                ), //i
    .io_passthrough (mac_4_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_0_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_129 mac_4_1 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_3_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_1_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_130 mac_4_2 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_3_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_2_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_131 mac_4_3 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_3_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_3_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_132 mac_4_4 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_3_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_4_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_133 mac_4_5 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_3_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_5_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_134 mac_4_6 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_3_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_6_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_135 mac_4_7 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_3_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_7_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_136 mac_4_8 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_3_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_8_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_137 mac_4_9 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_3_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_9_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_138 mac_4_10 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_3_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_4_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_10_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_139 mac_4_11 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_3_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_11_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_140 mac_4_12 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_3_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_12_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_141 mac_4_13 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_3_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_13_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_142 mac_4_14 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_3_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_14_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_143 mac_4_15 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_3_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_15_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_144 mac_4_16 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_3_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_16_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_145 mac_4_17 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_3_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_17_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_146 mac_4_18 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_3_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_18_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_147 mac_4_19 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_3_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_19_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_148 mac_4_20 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_3_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_20_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_149 mac_4_21 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_3_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_21_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_150 mac_4_22 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_3_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_22_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_151 mac_4_23 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_3_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_23_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_152 mac_4_24 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_3_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_24_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_153 mac_4_25 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_3_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_25_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_154 mac_4_26 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_3_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_26_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_155 mac_4_27 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_3_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_27_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_156 mac_4_28 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_3_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_28_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_157 mac_4_29 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_3_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_29_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_158 mac_4_30 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_3_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_30_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_159 mac_4_31 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_3_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_4_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_4_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_4_31_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_160 mac_5_0 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_4_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_5[7:0]                ), //i
    .io_passthrough (mac_5_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_0_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_161 mac_5_1 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_4_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_1_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_162 mac_5_2 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_4_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_2_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_163 mac_5_3 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_4_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_3_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_164 mac_5_4 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_4_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_4_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_165 mac_5_5 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_4_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_5_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_166 mac_5_6 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_4_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_6_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_167 mac_5_7 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_4_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_7_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_168 mac_5_8 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_4_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_8_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_169 mac_5_9 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_4_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_9_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_170 mac_5_10 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_4_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_5_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_10_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_171 mac_5_11 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_4_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_11_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_172 mac_5_12 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_4_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_12_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_173 mac_5_13 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_4_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_13_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_174 mac_5_14 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_4_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_14_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_175 mac_5_15 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_4_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_15_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_176 mac_5_16 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_4_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_16_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_177 mac_5_17 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_4_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_17_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_178 mac_5_18 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_4_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_18_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_179 mac_5_19 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_4_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_19_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_180 mac_5_20 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_4_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_20_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_181 mac_5_21 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_4_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_21_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_182 mac_5_22 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_4_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_22_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_183 mac_5_23 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_4_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_23_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_184 mac_5_24 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_4_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_24_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_185 mac_5_25 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_4_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_25_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_186 mac_5_26 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_4_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_26_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_187 mac_5_27 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_4_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_27_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_188 mac_5_28 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_4_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_28_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_189 mac_5_29 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_4_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_29_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_190 mac_5_30 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_4_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_30_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_191 mac_5_31 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_4_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_5_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_5_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_5_31_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_192 mac_6_0 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_5_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_6[7:0]                ), //i
    .io_passthrough (mac_6_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_0_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_193 mac_6_1 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_5_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_1_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_194 mac_6_2 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_5_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_2_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_195 mac_6_3 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_5_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_3_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_196 mac_6_4 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_5_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_4_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_197 mac_6_5 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_5_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_5_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_198 mac_6_6 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_5_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_6_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_199 mac_6_7 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_5_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_7_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_200 mac_6_8 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_5_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_8_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_201 mac_6_9 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_5_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_9_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_202 mac_6_10 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_5_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_6_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_10_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_203 mac_6_11 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_5_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_11_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_204 mac_6_12 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_5_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_12_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_205 mac_6_13 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_5_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_13_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_206 mac_6_14 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_5_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_14_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_207 mac_6_15 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_5_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_15_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_208 mac_6_16 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_5_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_16_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_209 mac_6_17 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_5_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_17_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_210 mac_6_18 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_5_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_18_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_211 mac_6_19 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_5_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_19_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_212 mac_6_20 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_5_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_20_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_213 mac_6_21 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_5_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_21_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_214 mac_6_22 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_5_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_22_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_215 mac_6_23 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_5_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_23_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_216 mac_6_24 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_5_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_24_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_217 mac_6_25 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_5_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_25_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_218 mac_6_26 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_5_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_26_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_219 mac_6_27 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_5_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_27_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_220 mac_6_28 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_5_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_28_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_221 mac_6_29 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_5_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_29_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_222 mac_6_30 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_5_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_30_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_223 mac_6_31 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_5_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_6_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_6_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_6_31_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_224 mac_7_0 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_6_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_7[7:0]                ), //i
    .io_passthrough (mac_7_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_0_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_225 mac_7_1 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_6_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_1_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_226 mac_7_2 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_6_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_2_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_227 mac_7_3 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_6_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_3_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_228 mac_7_4 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_6_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_4_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_229 mac_7_5 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_6_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_5_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_230 mac_7_6 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_6_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_6_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_231 mac_7_7 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_6_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_7_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_232 mac_7_8 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_6_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_8_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_233 mac_7_9 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_6_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_9_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_234 mac_7_10 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_6_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_7_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_10_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_235 mac_7_11 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_6_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_11_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_236 mac_7_12 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_6_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_12_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_237 mac_7_13 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_6_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_13_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_238 mac_7_14 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_6_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_14_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_239 mac_7_15 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_6_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_15_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_240 mac_7_16 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_6_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_16_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_241 mac_7_17 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_6_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_17_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_242 mac_7_18 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_6_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_18_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_243 mac_7_19 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_6_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_19_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_244 mac_7_20 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_6_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_20_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_245 mac_7_21 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_6_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_21_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_246 mac_7_22 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_6_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_22_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_247 mac_7_23 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_6_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_23_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_248 mac_7_24 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_6_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_24_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_249 mac_7_25 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_6_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_25_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_250 mac_7_26 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_6_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_26_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_251 mac_7_27 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_6_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_27_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_252 mac_7_28 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_6_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_28_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_253 mac_7_29 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_6_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_29_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_254 mac_7_30 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_6_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_30_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_255 mac_7_31 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_6_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_7_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_7_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_7_31_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_256 mac_8_0 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_7_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_8[7:0]                ), //i
    .io_passthrough (mac_8_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_0_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_257 mac_8_1 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_7_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_1_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_258 mac_8_2 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_7_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_2_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_259 mac_8_3 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_7_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_3_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_260 mac_8_4 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_7_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_4_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_261 mac_8_5 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_7_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_5_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_262 mac_8_6 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_7_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_6_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_263 mac_8_7 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_7_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_7_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_264 mac_8_8 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_7_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_8_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_265 mac_8_9 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_7_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_9_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_266 mac_8_10 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_7_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_8_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_10_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_267 mac_8_11 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_7_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_11_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_268 mac_8_12 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_7_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_12_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_269 mac_8_13 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_7_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_13_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_270 mac_8_14 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_7_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_14_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_271 mac_8_15 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_7_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_15_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_272 mac_8_16 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_7_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_16_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_273 mac_8_17 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_7_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_17_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_274 mac_8_18 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_7_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_18_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_275 mac_8_19 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_7_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_19_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_276 mac_8_20 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_7_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_20_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_277 mac_8_21 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_7_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_21_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_278 mac_8_22 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_7_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_22_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_279 mac_8_23 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_7_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_23_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_280 mac_8_24 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_7_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_24_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_281 mac_8_25 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_7_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_25_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_282 mac_8_26 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_7_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_26_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_283 mac_8_27 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_7_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_27_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_284 mac_8_28 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_7_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_28_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_285 mac_8_29 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_7_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_29_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_286 mac_8_30 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_7_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_30_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_287 mac_8_31 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_7_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_8_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_8_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_8_31_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_288 mac_9_0 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_8_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_9[7:0]                ), //i
    .io_passthrough (mac_9_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_0_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_289 mac_9_1 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_8_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_1_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_290 mac_9_2 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_8_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_2_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_291 mac_9_3 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_8_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_3_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_292 mac_9_4 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_8_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_4_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_293 mac_9_5 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_8_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_5_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_294 mac_9_6 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_8_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_6_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_295 mac_9_7 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_8_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_7_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_296 mac_9_8 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_8_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_8_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_297 mac_9_9 (
    .io_load        (io_load                    ), //i
    .io_mulInput    (mac_8_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_9_io_macOut[7:0]     ), //o
    .clk            (clk                        ), //i
    .reset          (reset                      )  //i
  );
  MAC_298 mac_9_10 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_8_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_9_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_10_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_299 mac_9_11 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_8_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_11_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_300 mac_9_12 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_8_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_12_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_301 mac_9_13 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_8_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_13_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_302 mac_9_14 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_8_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_14_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_303 mac_9_15 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_8_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_15_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_304 mac_9_16 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_8_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_16_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_305 mac_9_17 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_8_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_17_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_306 mac_9_18 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_8_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_18_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_307 mac_9_19 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_8_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_19_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_308 mac_9_20 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_8_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_20_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_309 mac_9_21 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_8_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_21_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_310 mac_9_22 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_8_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_22_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_311 mac_9_23 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_8_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_23_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_312 mac_9_24 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_8_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_24_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_313 mac_9_25 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_8_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_25_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_314 mac_9_26 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_8_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_26_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_315 mac_9_27 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_8_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_27_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_316 mac_9_28 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_8_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_28_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_317 mac_9_29 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_8_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_29_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_318 mac_9_30 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_8_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_30_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_319 mac_9_31 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_8_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_9_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_9_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_9_31_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_320 mac_10_0 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_9_0_io_passthrough[7:0] ), //i
    .io_addInput    (bias_10[7:0]                ), //i
    .io_passthrough (mac_10_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_0_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_321 mac_10_1 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_9_1_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_1_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_322 mac_10_2 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_9_2_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_2_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_323 mac_10_3 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_9_3_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_3_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_324 mac_10_4 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_9_4_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_4_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_325 mac_10_5 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_9_5_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_5_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_326 mac_10_6 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_9_6_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_6_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_327 mac_10_7 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_9_7_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_7_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_328 mac_10_8 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_9_8_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_8_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_329 mac_10_9 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_9_9_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_9_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_330 mac_10_10 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_9_10_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_10_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_10_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_331 mac_10_11 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_9_11_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_11_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_332 mac_10_12 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_9_12_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_12_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_333 mac_10_13 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_9_13_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_13_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_334 mac_10_14 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_9_14_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_14_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_335 mac_10_15 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_9_15_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_15_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_336 mac_10_16 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_9_16_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_16_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_337 mac_10_17 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_9_17_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_17_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_338 mac_10_18 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_9_18_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_18_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_339 mac_10_19 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_9_19_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_19_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_340 mac_10_20 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_9_20_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_20_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_341 mac_10_21 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_9_21_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_21_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_342 mac_10_22 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_9_22_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_22_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_343 mac_10_23 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_9_23_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_23_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_344 mac_10_24 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_9_24_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_24_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_345 mac_10_25 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_9_25_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_25_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_346 mac_10_26 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_9_26_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_26_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_347 mac_10_27 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_9_27_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_27_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_348 mac_10_28 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_9_28_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_28_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_349 mac_10_29 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_9_29_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_29_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_350 mac_10_30 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_9_30_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_30_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_351 mac_10_31 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_9_31_io_passthrough[7:0] ), //i
    .io_addInput    (mac_10_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_10_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_10_31_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_352 mac_11_0 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_10_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_11[7:0]                ), //i
    .io_passthrough (mac_11_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_0_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_353 mac_11_1 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_10_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_1_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_354 mac_11_2 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_10_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_2_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_355 mac_11_3 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_10_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_3_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_356 mac_11_4 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_10_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_4_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_357 mac_11_5 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_10_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_5_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_358 mac_11_6 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_10_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_6_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_359 mac_11_7 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_10_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_7_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_360 mac_11_8 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_10_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_8_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_361 mac_11_9 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_10_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_9_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_362 mac_11_10 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_10_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_11_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_10_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_363 mac_11_11 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_10_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_11_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_364 mac_11_12 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_10_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_12_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_365 mac_11_13 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_10_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_13_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_366 mac_11_14 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_10_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_14_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_367 mac_11_15 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_10_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_15_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_368 mac_11_16 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_10_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_16_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_369 mac_11_17 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_10_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_17_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_370 mac_11_18 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_10_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_18_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_371 mac_11_19 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_10_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_19_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_372 mac_11_20 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_10_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_20_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_373 mac_11_21 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_10_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_21_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_374 mac_11_22 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_10_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_22_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_375 mac_11_23 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_10_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_23_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_376 mac_11_24 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_10_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_24_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_377 mac_11_25 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_10_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_25_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_378 mac_11_26 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_10_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_26_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_379 mac_11_27 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_10_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_27_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_380 mac_11_28 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_10_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_28_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_381 mac_11_29 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_10_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_29_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_382 mac_11_30 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_10_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_30_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_383 mac_11_31 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_10_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_11_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_11_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_11_31_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_384 mac_12_0 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_11_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_12[7:0]                ), //i
    .io_passthrough (mac_12_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_0_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_385 mac_12_1 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_11_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_1_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_386 mac_12_2 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_11_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_2_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_387 mac_12_3 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_11_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_3_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_388 mac_12_4 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_11_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_4_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_389 mac_12_5 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_11_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_5_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_390 mac_12_6 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_11_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_6_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_391 mac_12_7 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_11_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_7_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_392 mac_12_8 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_11_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_8_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_393 mac_12_9 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_11_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_9_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_394 mac_12_10 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_11_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_12_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_10_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_395 mac_12_11 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_11_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_11_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_396 mac_12_12 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_11_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_12_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_397 mac_12_13 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_11_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_13_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_398 mac_12_14 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_11_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_14_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_399 mac_12_15 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_11_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_15_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_400 mac_12_16 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_11_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_16_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_401 mac_12_17 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_11_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_17_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_402 mac_12_18 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_11_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_18_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_403 mac_12_19 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_11_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_19_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_404 mac_12_20 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_11_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_20_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_405 mac_12_21 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_11_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_21_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_406 mac_12_22 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_11_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_22_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_407 mac_12_23 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_11_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_23_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_408 mac_12_24 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_11_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_24_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_409 mac_12_25 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_11_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_25_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_410 mac_12_26 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_11_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_26_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_411 mac_12_27 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_11_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_27_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_412 mac_12_28 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_11_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_28_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_413 mac_12_29 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_11_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_29_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_414 mac_12_30 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_11_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_30_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_415 mac_12_31 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_11_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_12_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_12_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_12_31_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_416 mac_13_0 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_12_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_13[7:0]                ), //i
    .io_passthrough (mac_13_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_0_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_417 mac_13_1 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_12_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_1_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_418 mac_13_2 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_12_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_2_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_419 mac_13_3 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_12_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_3_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_420 mac_13_4 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_12_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_4_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_421 mac_13_5 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_12_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_5_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_422 mac_13_6 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_12_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_6_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_423 mac_13_7 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_12_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_7_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_424 mac_13_8 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_12_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_8_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_425 mac_13_9 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_12_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_9_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_426 mac_13_10 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_12_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_13_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_10_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_427 mac_13_11 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_12_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_11_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_428 mac_13_12 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_12_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_12_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_429 mac_13_13 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_12_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_13_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_430 mac_13_14 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_12_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_14_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_431 mac_13_15 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_12_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_15_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_432 mac_13_16 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_12_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_16_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_433 mac_13_17 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_12_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_17_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_434 mac_13_18 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_12_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_18_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_435 mac_13_19 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_12_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_19_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_436 mac_13_20 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_12_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_20_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_437 mac_13_21 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_12_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_21_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_438 mac_13_22 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_12_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_22_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_439 mac_13_23 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_12_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_23_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_440 mac_13_24 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_12_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_24_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_441 mac_13_25 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_12_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_25_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_442 mac_13_26 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_12_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_26_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_443 mac_13_27 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_12_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_27_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_444 mac_13_28 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_12_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_28_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_445 mac_13_29 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_12_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_29_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_446 mac_13_30 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_12_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_30_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_447 mac_13_31 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_12_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_13_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_13_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_13_31_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_448 mac_14_0 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_13_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_14[7:0]                ), //i
    .io_passthrough (mac_14_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_0_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_449 mac_14_1 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_13_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_1_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_450 mac_14_2 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_13_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_2_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_451 mac_14_3 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_13_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_3_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_452 mac_14_4 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_13_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_4_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_453 mac_14_5 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_13_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_5_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_454 mac_14_6 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_13_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_6_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_455 mac_14_7 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_13_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_7_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_456 mac_14_8 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_13_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_8_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_457 mac_14_9 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_13_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_9_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_458 mac_14_10 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_13_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_14_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_10_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_459 mac_14_11 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_13_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_11_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_460 mac_14_12 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_13_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_12_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_461 mac_14_13 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_13_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_13_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_462 mac_14_14 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_13_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_14_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_463 mac_14_15 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_13_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_15_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_464 mac_14_16 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_13_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_16_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_465 mac_14_17 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_13_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_17_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_466 mac_14_18 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_13_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_18_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_467 mac_14_19 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_13_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_19_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_468 mac_14_20 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_13_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_20_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_469 mac_14_21 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_13_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_21_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_470 mac_14_22 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_13_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_22_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_471 mac_14_23 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_13_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_23_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_472 mac_14_24 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_13_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_24_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_473 mac_14_25 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_13_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_25_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_474 mac_14_26 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_13_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_26_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_475 mac_14_27 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_13_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_27_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_476 mac_14_28 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_13_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_28_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_477 mac_14_29 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_13_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_29_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_478 mac_14_30 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_13_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_30_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_479 mac_14_31 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_13_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_14_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_14_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_14_31_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_480 mac_15_0 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_14_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_15[7:0]                ), //i
    .io_passthrough (mac_15_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_0_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_481 mac_15_1 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_14_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_1_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_482 mac_15_2 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_14_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_2_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_483 mac_15_3 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_14_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_3_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_484 mac_15_4 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_14_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_4_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_485 mac_15_5 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_14_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_5_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_486 mac_15_6 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_14_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_6_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_487 mac_15_7 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_14_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_7_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_488 mac_15_8 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_14_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_8_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_489 mac_15_9 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_14_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_9_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_490 mac_15_10 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_14_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_15_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_10_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_491 mac_15_11 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_14_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_11_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_492 mac_15_12 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_14_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_12_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_493 mac_15_13 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_14_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_13_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_494 mac_15_14 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_14_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_14_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_495 mac_15_15 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_14_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_15_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_496 mac_15_16 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_14_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_16_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_497 mac_15_17 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_14_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_17_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_498 mac_15_18 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_14_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_18_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_499 mac_15_19 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_14_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_19_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_500 mac_15_20 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_14_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_20_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_501 mac_15_21 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_14_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_21_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_502 mac_15_22 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_14_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_22_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_503 mac_15_23 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_14_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_23_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_504 mac_15_24 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_14_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_24_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_505 mac_15_25 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_14_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_25_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_506 mac_15_26 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_14_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_26_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_507 mac_15_27 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_14_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_27_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_508 mac_15_28 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_14_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_28_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_509 mac_15_29 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_14_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_29_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_510 mac_15_30 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_14_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_30_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_511 mac_15_31 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_14_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_15_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_15_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_15_31_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_512 mac_16_0 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_15_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_16[7:0]                ), //i
    .io_passthrough (mac_16_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_0_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_513 mac_16_1 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_15_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_1_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_514 mac_16_2 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_15_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_2_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_515 mac_16_3 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_15_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_3_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_516 mac_16_4 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_15_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_4_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_517 mac_16_5 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_15_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_5_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_518 mac_16_6 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_15_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_6_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_519 mac_16_7 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_15_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_7_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_520 mac_16_8 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_15_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_8_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_521 mac_16_9 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_15_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_9_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_522 mac_16_10 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_15_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_16_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_10_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_523 mac_16_11 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_15_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_11_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_524 mac_16_12 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_15_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_12_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_525 mac_16_13 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_15_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_13_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_526 mac_16_14 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_15_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_14_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_527 mac_16_15 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_15_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_15_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_528 mac_16_16 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_15_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_16_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_529 mac_16_17 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_15_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_17_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_530 mac_16_18 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_15_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_18_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_531 mac_16_19 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_15_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_19_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_532 mac_16_20 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_15_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_20_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_533 mac_16_21 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_15_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_21_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_534 mac_16_22 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_15_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_22_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_535 mac_16_23 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_15_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_23_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_536 mac_16_24 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_15_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_24_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_537 mac_16_25 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_15_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_25_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_538 mac_16_26 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_15_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_26_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_539 mac_16_27 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_15_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_27_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_540 mac_16_28 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_15_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_28_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_541 mac_16_29 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_15_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_29_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_542 mac_16_30 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_15_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_30_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_543 mac_16_31 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_15_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_16_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_16_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_16_31_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_544 mac_17_0 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_16_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_17[7:0]                ), //i
    .io_passthrough (mac_17_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_0_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_545 mac_17_1 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_16_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_1_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_546 mac_17_2 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_16_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_2_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_547 mac_17_3 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_16_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_3_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_548 mac_17_4 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_16_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_4_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_549 mac_17_5 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_16_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_5_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_550 mac_17_6 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_16_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_6_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_551 mac_17_7 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_16_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_7_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_552 mac_17_8 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_16_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_8_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_553 mac_17_9 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_16_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_9_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_554 mac_17_10 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_16_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_17_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_10_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_555 mac_17_11 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_16_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_11_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_556 mac_17_12 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_16_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_12_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_557 mac_17_13 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_16_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_13_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_558 mac_17_14 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_16_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_14_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_559 mac_17_15 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_16_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_15_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_560 mac_17_16 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_16_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_16_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_561 mac_17_17 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_16_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_17_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_562 mac_17_18 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_16_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_18_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_563 mac_17_19 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_16_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_19_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_564 mac_17_20 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_16_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_20_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_565 mac_17_21 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_16_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_21_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_566 mac_17_22 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_16_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_22_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_567 mac_17_23 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_16_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_23_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_568 mac_17_24 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_16_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_24_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_569 mac_17_25 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_16_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_25_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_570 mac_17_26 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_16_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_26_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_571 mac_17_27 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_16_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_27_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_572 mac_17_28 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_16_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_28_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_573 mac_17_29 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_16_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_29_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_574 mac_17_30 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_16_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_30_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_575 mac_17_31 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_16_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_17_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_17_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_17_31_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_576 mac_18_0 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_17_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_18[7:0]                ), //i
    .io_passthrough (mac_18_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_0_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_577 mac_18_1 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_17_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_1_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_578 mac_18_2 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_17_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_2_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_579 mac_18_3 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_17_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_3_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_580 mac_18_4 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_17_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_4_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_581 mac_18_5 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_17_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_5_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_582 mac_18_6 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_17_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_6_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_583 mac_18_7 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_17_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_7_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_584 mac_18_8 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_17_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_8_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_585 mac_18_9 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_17_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_9_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_586 mac_18_10 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_17_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_18_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_10_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_587 mac_18_11 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_17_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_11_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_588 mac_18_12 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_17_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_12_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_589 mac_18_13 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_17_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_13_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_590 mac_18_14 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_17_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_14_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_591 mac_18_15 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_17_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_15_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_592 mac_18_16 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_17_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_16_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_593 mac_18_17 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_17_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_17_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_594 mac_18_18 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_17_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_18_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_595 mac_18_19 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_17_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_19_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_596 mac_18_20 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_17_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_20_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_597 mac_18_21 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_17_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_21_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_598 mac_18_22 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_17_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_22_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_599 mac_18_23 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_17_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_23_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_600 mac_18_24 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_17_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_24_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_601 mac_18_25 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_17_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_25_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_602 mac_18_26 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_17_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_26_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_603 mac_18_27 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_17_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_27_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_604 mac_18_28 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_17_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_28_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_605 mac_18_29 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_17_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_29_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_606 mac_18_30 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_17_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_30_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_607 mac_18_31 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_17_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_18_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_18_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_18_31_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_608 mac_19_0 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_18_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_19[7:0]                ), //i
    .io_passthrough (mac_19_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_0_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_609 mac_19_1 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_18_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_1_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_610 mac_19_2 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_18_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_2_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_611 mac_19_3 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_18_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_3_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_612 mac_19_4 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_18_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_4_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_613 mac_19_5 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_18_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_5_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_614 mac_19_6 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_18_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_6_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_615 mac_19_7 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_18_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_7_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_616 mac_19_8 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_18_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_8_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_617 mac_19_9 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_18_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_9_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_618 mac_19_10 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_18_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_19_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_10_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_619 mac_19_11 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_18_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_11_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_620 mac_19_12 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_18_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_12_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_621 mac_19_13 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_18_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_13_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_622 mac_19_14 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_18_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_14_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_623 mac_19_15 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_18_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_15_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_624 mac_19_16 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_18_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_16_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_625 mac_19_17 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_18_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_17_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_626 mac_19_18 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_18_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_18_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_627 mac_19_19 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_18_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_19_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_628 mac_19_20 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_18_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_20_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_629 mac_19_21 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_18_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_21_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_630 mac_19_22 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_18_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_22_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_631 mac_19_23 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_18_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_23_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_632 mac_19_24 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_18_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_24_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_633 mac_19_25 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_18_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_25_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_634 mac_19_26 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_18_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_26_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_635 mac_19_27 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_18_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_27_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_636 mac_19_28 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_18_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_28_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_637 mac_19_29 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_18_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_29_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_638 mac_19_30 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_18_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_30_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_639 mac_19_31 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_18_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_19_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_19_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_19_31_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_640 mac_20_0 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_19_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_20[7:0]                ), //i
    .io_passthrough (mac_20_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_0_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_641 mac_20_1 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_19_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_1_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_642 mac_20_2 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_19_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_2_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_643 mac_20_3 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_19_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_3_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_644 mac_20_4 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_19_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_4_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_645 mac_20_5 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_19_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_5_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_646 mac_20_6 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_19_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_6_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_647 mac_20_7 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_19_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_7_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_648 mac_20_8 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_19_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_8_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_649 mac_20_9 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_19_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_9_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_650 mac_20_10 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_19_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_20_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_10_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_651 mac_20_11 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_19_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_11_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_652 mac_20_12 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_19_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_12_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_653 mac_20_13 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_19_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_13_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_654 mac_20_14 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_19_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_14_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_655 mac_20_15 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_19_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_15_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_656 mac_20_16 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_19_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_16_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_657 mac_20_17 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_19_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_17_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_658 mac_20_18 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_19_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_18_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_659 mac_20_19 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_19_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_19_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_660 mac_20_20 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_19_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_20_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_661 mac_20_21 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_19_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_21_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_662 mac_20_22 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_19_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_22_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_663 mac_20_23 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_19_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_23_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_664 mac_20_24 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_19_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_24_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_665 mac_20_25 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_19_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_25_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_666 mac_20_26 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_19_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_26_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_667 mac_20_27 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_19_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_27_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_668 mac_20_28 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_19_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_28_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_669 mac_20_29 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_19_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_29_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_670 mac_20_30 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_19_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_30_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_671 mac_20_31 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_19_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_20_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_20_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_20_31_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_672 mac_21_0 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_20_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_21[7:0]                ), //i
    .io_passthrough (mac_21_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_0_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_673 mac_21_1 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_20_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_1_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_674 mac_21_2 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_20_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_2_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_675 mac_21_3 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_20_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_3_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_676 mac_21_4 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_20_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_4_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_677 mac_21_5 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_20_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_5_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_678 mac_21_6 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_20_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_6_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_679 mac_21_7 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_20_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_7_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_680 mac_21_8 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_20_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_8_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_681 mac_21_9 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_20_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_9_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_682 mac_21_10 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_20_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_21_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_10_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_683 mac_21_11 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_20_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_11_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_684 mac_21_12 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_20_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_12_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_685 mac_21_13 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_20_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_13_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_686 mac_21_14 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_20_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_14_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_687 mac_21_15 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_20_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_15_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_688 mac_21_16 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_20_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_16_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_689 mac_21_17 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_20_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_17_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_690 mac_21_18 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_20_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_18_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_691 mac_21_19 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_20_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_19_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_692 mac_21_20 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_20_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_20_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_693 mac_21_21 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_20_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_21_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_694 mac_21_22 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_20_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_22_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_695 mac_21_23 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_20_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_23_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_696 mac_21_24 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_20_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_24_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_697 mac_21_25 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_20_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_25_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_698 mac_21_26 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_20_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_26_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_699 mac_21_27 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_20_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_27_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_700 mac_21_28 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_20_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_28_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_701 mac_21_29 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_20_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_29_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_702 mac_21_30 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_20_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_30_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_703 mac_21_31 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_20_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_21_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_21_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_21_31_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_704 mac_22_0 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_21_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_22[7:0]                ), //i
    .io_passthrough (mac_22_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_0_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_705 mac_22_1 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_21_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_1_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_706 mac_22_2 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_21_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_2_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_707 mac_22_3 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_21_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_3_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_708 mac_22_4 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_21_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_4_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_709 mac_22_5 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_21_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_5_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_710 mac_22_6 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_21_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_6_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_711 mac_22_7 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_21_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_7_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_712 mac_22_8 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_21_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_8_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_713 mac_22_9 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_21_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_9_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_714 mac_22_10 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_21_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_22_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_10_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_715 mac_22_11 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_21_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_11_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_716 mac_22_12 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_21_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_12_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_717 mac_22_13 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_21_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_13_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_718 mac_22_14 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_21_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_14_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_719 mac_22_15 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_21_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_15_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_720 mac_22_16 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_21_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_16_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_721 mac_22_17 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_21_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_17_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_722 mac_22_18 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_21_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_18_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_723 mac_22_19 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_21_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_19_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_724 mac_22_20 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_21_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_20_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_725 mac_22_21 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_21_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_21_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_726 mac_22_22 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_21_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_22_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_727 mac_22_23 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_21_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_23_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_728 mac_22_24 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_21_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_24_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_729 mac_22_25 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_21_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_25_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_730 mac_22_26 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_21_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_26_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_731 mac_22_27 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_21_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_27_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_732 mac_22_28 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_21_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_28_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_733 mac_22_29 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_21_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_29_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_734 mac_22_30 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_21_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_30_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_735 mac_22_31 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_21_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_22_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_22_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_22_31_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_736 mac_23_0 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_22_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_23[7:0]                ), //i
    .io_passthrough (mac_23_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_0_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_737 mac_23_1 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_22_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_1_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_738 mac_23_2 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_22_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_2_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_739 mac_23_3 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_22_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_3_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_740 mac_23_4 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_22_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_4_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_741 mac_23_5 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_22_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_5_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_742 mac_23_6 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_22_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_6_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_743 mac_23_7 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_22_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_7_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_744 mac_23_8 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_22_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_8_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_745 mac_23_9 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_22_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_9_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_746 mac_23_10 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_22_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_23_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_10_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_747 mac_23_11 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_22_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_11_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_748 mac_23_12 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_22_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_12_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_749 mac_23_13 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_22_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_13_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_750 mac_23_14 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_22_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_14_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_751 mac_23_15 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_22_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_15_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_752 mac_23_16 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_22_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_16_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_753 mac_23_17 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_22_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_17_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_754 mac_23_18 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_22_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_18_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_755 mac_23_19 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_22_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_19_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_756 mac_23_20 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_22_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_20_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_757 mac_23_21 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_22_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_21_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_758 mac_23_22 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_22_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_22_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_759 mac_23_23 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_22_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_23_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_760 mac_23_24 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_22_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_24_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_761 mac_23_25 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_22_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_25_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_762 mac_23_26 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_22_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_26_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_763 mac_23_27 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_22_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_27_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_764 mac_23_28 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_22_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_28_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_765 mac_23_29 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_22_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_29_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_766 mac_23_30 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_22_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_30_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_767 mac_23_31 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_22_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_23_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_23_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_23_31_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_768 mac_24_0 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_23_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_24[7:0]                ), //i
    .io_passthrough (mac_24_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_0_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_769 mac_24_1 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_23_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_1_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_770 mac_24_2 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_23_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_2_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_771 mac_24_3 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_23_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_3_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_772 mac_24_4 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_23_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_4_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_773 mac_24_5 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_23_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_5_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_774 mac_24_6 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_23_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_6_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_775 mac_24_7 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_23_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_7_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_776 mac_24_8 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_23_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_8_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_777 mac_24_9 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_23_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_9_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_778 mac_24_10 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_23_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_24_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_10_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_779 mac_24_11 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_23_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_11_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_780 mac_24_12 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_23_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_12_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_781 mac_24_13 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_23_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_13_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_782 mac_24_14 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_23_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_14_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_783 mac_24_15 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_23_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_15_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_784 mac_24_16 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_23_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_16_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_785 mac_24_17 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_23_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_17_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_786 mac_24_18 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_23_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_18_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_787 mac_24_19 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_23_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_19_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_788 mac_24_20 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_23_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_20_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_789 mac_24_21 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_23_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_21_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_790 mac_24_22 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_23_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_22_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_791 mac_24_23 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_23_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_23_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_792 mac_24_24 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_23_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_24_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_793 mac_24_25 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_23_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_25_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_794 mac_24_26 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_23_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_26_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_795 mac_24_27 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_23_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_27_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_796 mac_24_28 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_23_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_28_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_797 mac_24_29 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_23_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_29_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_798 mac_24_30 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_23_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_30_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_799 mac_24_31 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_23_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_24_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_24_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_24_31_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_800 mac_25_0 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_24_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_25[7:0]                ), //i
    .io_passthrough (mac_25_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_0_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_801 mac_25_1 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_24_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_1_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_802 mac_25_2 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_24_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_2_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_803 mac_25_3 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_24_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_3_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_804 mac_25_4 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_24_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_4_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_805 mac_25_5 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_24_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_5_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_806 mac_25_6 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_24_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_6_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_807 mac_25_7 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_24_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_7_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_808 mac_25_8 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_24_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_8_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_809 mac_25_9 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_24_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_9_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_810 mac_25_10 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_24_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_25_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_10_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_811 mac_25_11 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_24_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_11_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_812 mac_25_12 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_24_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_12_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_813 mac_25_13 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_24_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_13_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_814 mac_25_14 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_24_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_14_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_815 mac_25_15 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_24_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_15_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_816 mac_25_16 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_24_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_16_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_817 mac_25_17 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_24_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_17_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_818 mac_25_18 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_24_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_18_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_819 mac_25_19 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_24_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_19_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_820 mac_25_20 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_24_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_20_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_821 mac_25_21 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_24_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_21_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_822 mac_25_22 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_24_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_22_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_823 mac_25_23 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_24_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_23_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_824 mac_25_24 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_24_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_24_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_825 mac_25_25 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_24_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_25_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_826 mac_25_26 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_24_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_26_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_827 mac_25_27 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_24_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_27_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_828 mac_25_28 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_24_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_28_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_829 mac_25_29 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_24_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_29_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_830 mac_25_30 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_24_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_30_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_831 mac_25_31 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_24_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_25_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_25_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_25_31_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_832 mac_26_0 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_25_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_26[7:0]                ), //i
    .io_passthrough (mac_26_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_0_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_833 mac_26_1 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_25_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_1_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_834 mac_26_2 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_25_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_2_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_835 mac_26_3 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_25_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_3_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_836 mac_26_4 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_25_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_4_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_837 mac_26_5 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_25_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_5_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_838 mac_26_6 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_25_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_6_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_839 mac_26_7 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_25_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_7_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_840 mac_26_8 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_25_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_8_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_841 mac_26_9 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_25_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_9_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_842 mac_26_10 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_25_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_26_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_10_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_843 mac_26_11 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_25_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_11_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_844 mac_26_12 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_25_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_12_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_845 mac_26_13 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_25_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_13_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_846 mac_26_14 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_25_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_14_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_847 mac_26_15 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_25_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_15_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_848 mac_26_16 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_25_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_16_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_849 mac_26_17 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_25_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_17_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_850 mac_26_18 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_25_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_18_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_851 mac_26_19 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_25_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_19_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_852 mac_26_20 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_25_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_20_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_853 mac_26_21 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_25_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_21_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_854 mac_26_22 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_25_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_22_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_855 mac_26_23 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_25_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_23_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_856 mac_26_24 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_25_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_24_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_857 mac_26_25 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_25_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_25_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_858 mac_26_26 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_25_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_26_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_859 mac_26_27 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_25_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_27_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_860 mac_26_28 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_25_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_28_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_861 mac_26_29 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_25_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_29_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_862 mac_26_30 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_25_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_30_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_863 mac_26_31 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_25_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_26_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_26_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_26_31_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_864 mac_27_0 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_26_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_27[7:0]                ), //i
    .io_passthrough (mac_27_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_0_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_865 mac_27_1 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_26_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_1_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_866 mac_27_2 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_26_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_2_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_867 mac_27_3 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_26_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_3_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_868 mac_27_4 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_26_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_4_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_869 mac_27_5 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_26_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_5_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_870 mac_27_6 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_26_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_6_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_871 mac_27_7 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_26_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_7_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_872 mac_27_8 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_26_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_8_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_873 mac_27_9 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_26_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_9_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_874 mac_27_10 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_26_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_27_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_10_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_875 mac_27_11 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_26_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_11_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_876 mac_27_12 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_26_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_12_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_877 mac_27_13 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_26_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_13_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_878 mac_27_14 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_26_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_14_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_879 mac_27_15 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_26_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_15_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_880 mac_27_16 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_26_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_16_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_881 mac_27_17 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_26_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_17_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_882 mac_27_18 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_26_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_18_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_883 mac_27_19 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_26_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_19_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_884 mac_27_20 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_26_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_20_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_885 mac_27_21 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_26_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_21_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_886 mac_27_22 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_26_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_22_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_887 mac_27_23 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_26_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_23_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_888 mac_27_24 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_26_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_24_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_889 mac_27_25 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_26_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_25_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_890 mac_27_26 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_26_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_26_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_891 mac_27_27 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_26_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_27_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_892 mac_27_28 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_26_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_28_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_893 mac_27_29 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_26_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_29_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_894 mac_27_30 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_26_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_30_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_895 mac_27_31 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_26_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_27_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_27_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_27_31_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_896 mac_28_0 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_27_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_28[7:0]                ), //i
    .io_passthrough (mac_28_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_0_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_897 mac_28_1 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_27_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_1_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_898 mac_28_2 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_27_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_2_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_899 mac_28_3 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_27_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_3_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_900 mac_28_4 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_27_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_4_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_901 mac_28_5 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_27_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_5_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_902 mac_28_6 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_27_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_6_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_903 mac_28_7 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_27_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_7_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_904 mac_28_8 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_27_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_8_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_905 mac_28_9 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_27_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_9_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_906 mac_28_10 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_27_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_28_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_10_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_907 mac_28_11 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_27_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_11_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_908 mac_28_12 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_27_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_12_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_909 mac_28_13 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_27_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_13_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_910 mac_28_14 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_27_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_14_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_911 mac_28_15 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_27_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_15_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_912 mac_28_16 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_27_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_16_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_913 mac_28_17 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_27_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_17_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_914 mac_28_18 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_27_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_18_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_915 mac_28_19 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_27_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_19_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_916 mac_28_20 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_27_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_20_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_917 mac_28_21 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_27_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_21_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_918 mac_28_22 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_27_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_22_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_919 mac_28_23 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_27_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_23_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_920 mac_28_24 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_27_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_24_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_921 mac_28_25 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_27_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_25_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_922 mac_28_26 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_27_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_26_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_923 mac_28_27 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_27_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_27_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_924 mac_28_28 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_27_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_28_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_925 mac_28_29 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_27_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_29_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_926 mac_28_30 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_27_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_30_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_927 mac_28_31 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_27_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_28_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_28_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_28_31_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_928 mac_29_0 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_28_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_29[7:0]                ), //i
    .io_passthrough (mac_29_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_0_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_929 mac_29_1 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_28_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_1_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_930 mac_29_2 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_28_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_2_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_931 mac_29_3 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_28_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_3_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_932 mac_29_4 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_28_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_4_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_933 mac_29_5 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_28_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_5_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_934 mac_29_6 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_28_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_6_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_935 mac_29_7 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_28_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_7_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_936 mac_29_8 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_28_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_8_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_937 mac_29_9 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_28_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_9_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_938 mac_29_10 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_28_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_29_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_10_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_939 mac_29_11 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_28_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_11_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_940 mac_29_12 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_28_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_12_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_941 mac_29_13 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_28_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_13_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_942 mac_29_14 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_28_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_14_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_943 mac_29_15 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_28_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_15_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_944 mac_29_16 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_28_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_16_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_945 mac_29_17 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_28_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_17_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_946 mac_29_18 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_28_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_18_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_947 mac_29_19 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_28_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_19_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_948 mac_29_20 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_28_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_20_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_949 mac_29_21 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_28_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_21_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_950 mac_29_22 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_28_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_22_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_951 mac_29_23 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_28_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_23_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_952 mac_29_24 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_28_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_24_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_953 mac_29_25 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_28_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_25_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_954 mac_29_26 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_28_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_26_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_955 mac_29_27 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_28_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_27_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_956 mac_29_28 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_28_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_28_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_957 mac_29_29 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_28_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_29_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_958 mac_29_30 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_28_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_30_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_959 mac_29_31 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_28_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_29_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_29_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_29_31_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_960 mac_30_0 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_29_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_30[7:0]                ), //i
    .io_passthrough (mac_30_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_0_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_961 mac_30_1 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_29_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_1_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_962 mac_30_2 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_29_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_2_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_963 mac_30_3 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_29_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_3_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_964 mac_30_4 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_29_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_4_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_965 mac_30_5 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_29_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_5_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_966 mac_30_6 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_29_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_6_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_967 mac_30_7 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_29_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_7_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_968 mac_30_8 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_29_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_8_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_969 mac_30_9 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_29_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_9_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_970 mac_30_10 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_29_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_30_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_10_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_971 mac_30_11 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_29_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_11_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_972 mac_30_12 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_29_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_12_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_973 mac_30_13 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_29_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_13_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_974 mac_30_14 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_29_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_14_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_975 mac_30_15 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_29_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_15_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_976 mac_30_16 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_29_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_16_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_977 mac_30_17 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_29_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_17_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_978 mac_30_18 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_29_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_18_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_979 mac_30_19 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_29_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_19_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_980 mac_30_20 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_29_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_20_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_981 mac_30_21 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_29_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_21_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_982 mac_30_22 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_29_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_22_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_983 mac_30_23 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_29_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_23_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_984 mac_30_24 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_29_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_24_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_985 mac_30_25 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_29_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_25_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_986 mac_30_26 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_29_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_26_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_987 mac_30_27 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_29_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_27_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_988 mac_30_28 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_29_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_28_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_989 mac_30_29 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_29_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_29_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_990 mac_30_30 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_29_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_30_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_991 mac_30_31 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_29_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_30_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_30_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_30_31_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_992 mac_31_0 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_30_0_io_passthrough[7:0]), //i
    .io_addInput    (bias_31[7:0]                ), //i
    .io_passthrough (mac_31_0_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_0_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_993 mac_31_1 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_30_1_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_0_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_1_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_1_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_994 mac_31_2 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_30_2_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_1_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_2_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_2_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_995 mac_31_3 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_30_3_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_2_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_3_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_3_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_996 mac_31_4 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_30_4_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_3_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_4_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_4_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_997 mac_31_5 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_30_5_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_4_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_5_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_5_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_998 mac_31_6 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_30_6_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_5_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_6_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_6_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_999 mac_31_7 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_30_7_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_6_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_7_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_7_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_1000 mac_31_8 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_30_8_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_7_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_8_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_8_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_1001 mac_31_9 (
    .io_load        (io_load                     ), //i
    .io_mulInput    (mac_30_9_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_8_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_9_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_9_io_macOut[7:0]     ), //o
    .clk            (clk                         ), //i
    .reset          (reset                       )  //i
  );
  MAC_1002 mac_31_10 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_30_10_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_9_io_macOut[7:0]      ), //i
    .io_passthrough (mac_31_10_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_10_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_1003 mac_31_11 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_30_11_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_10_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_11_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_11_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_1004 mac_31_12 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_30_12_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_11_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_12_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_12_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_1005 mac_31_13 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_30_13_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_12_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_13_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_13_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_1006 mac_31_14 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_30_14_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_13_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_14_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_14_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_1007 mac_31_15 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_30_15_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_14_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_15_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_15_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_1008 mac_31_16 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_30_16_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_15_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_16_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_16_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_1009 mac_31_17 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_30_17_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_16_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_17_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_17_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_1010 mac_31_18 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_30_18_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_17_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_18_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_18_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_1011 mac_31_19 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_30_19_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_18_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_19_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_19_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_1012 mac_31_20 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_30_20_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_19_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_20_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_20_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_1013 mac_31_21 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_30_21_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_20_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_21_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_21_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_1014 mac_31_22 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_30_22_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_21_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_22_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_22_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_1015 mac_31_23 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_30_23_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_22_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_23_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_23_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_1016 mac_31_24 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_30_24_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_23_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_24_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_24_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_1017 mac_31_25 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_30_25_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_24_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_25_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_25_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_1018 mac_31_26 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_30_26_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_25_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_26_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_26_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_1019 mac_31_27 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_30_27_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_26_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_27_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_27_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_1020 mac_31_28 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_30_28_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_27_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_28_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_28_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_1021 mac_31_29 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_30_29_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_28_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_29_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_29_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_1022 mac_31_30 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_30_30_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_29_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_30_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_30_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  MAC_1023 mac_31_31 (
    .io_load        (io_load                      ), //i
    .io_mulInput    (mac_30_31_io_passthrough[7:0]), //i
    .io_addInput    (mac_31_30_io_macOut[7:0]     ), //i
    .io_passthrough (mac_31_31_io_passthrough[7:0]), //o
    .io_macOut      (mac_31_31_io_macOut[7:0]     ), //o
    .clk            (clk                          ), //i
    .reset          (reset                        )  //i
  );
  assign io_output_0 = toplevel_mac_0_31_io_macOut_delay_31;
  assign io_output_1 = toplevel_mac_1_31_io_macOut_delay_30;
  assign io_output_2 = toplevel_mac_2_31_io_macOut_delay_29;
  assign io_output_3 = toplevel_mac_3_31_io_macOut_delay_28;
  assign io_output_4 = toplevel_mac_4_31_io_macOut_delay_27;
  assign io_output_5 = toplevel_mac_5_31_io_macOut_delay_26;
  assign io_output_6 = toplevel_mac_6_31_io_macOut_delay_25;
  assign io_output_7 = toplevel_mac_7_31_io_macOut_delay_24;
  assign io_output_8 = toplevel_mac_8_31_io_macOut_delay_23;
  assign io_output_9 = toplevel_mac_9_31_io_macOut_delay_22;
  assign io_output_10 = toplevel_mac_10_31_io_macOut_delay_21;
  assign io_output_11 = toplevel_mac_11_31_io_macOut_delay_20;
  assign io_output_12 = toplevel_mac_12_31_io_macOut_delay_19;
  assign io_output_13 = toplevel_mac_13_31_io_macOut_delay_18;
  assign io_output_14 = toplevel_mac_14_31_io_macOut_delay_17;
  assign io_output_15 = toplevel_mac_15_31_io_macOut_delay_16;
  assign io_output_16 = toplevel_mac_16_31_io_macOut_delay_15;
  assign io_output_17 = toplevel_mac_17_31_io_macOut_delay_14;
  assign io_output_18 = toplevel_mac_18_31_io_macOut_delay_13;
  assign io_output_19 = toplevel_mac_19_31_io_macOut_delay_12;
  assign io_output_20 = toplevel_mac_20_31_io_macOut_delay_11;
  assign io_output_21 = toplevel_mac_21_31_io_macOut_delay_10;
  assign io_output_22 = toplevel_mac_22_31_io_macOut_delay_9;
  assign io_output_23 = toplevel_mac_23_31_io_macOut_delay_8;
  assign io_output_24 = toplevel_mac_24_31_io_macOut_delay_7;
  assign io_output_25 = toplevel_mac_25_31_io_macOut_delay_6;
  assign io_output_26 = toplevel_mac_26_31_io_macOut_delay_5;
  assign io_output_27 = toplevel_mac_27_31_io_macOut_delay_4;
  assign io_output_28 = toplevel_mac_28_31_io_macOut_delay_3;
  assign io_output_29 = toplevel_mac_29_31_io_macOut_delay_2;
  assign io_output_30 = toplevel_mac_30_31_io_macOut_delay_1;
  assign io_output_31 = mac_31_31_io_macOut;
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      bias_0 <= 8'h00;
      bias_1 <= 8'h00;
      bias_2 <= 8'h00;
      bias_3 <= 8'h00;
      bias_4 <= 8'h00;
      bias_5 <= 8'h00;
      bias_6 <= 8'h00;
      bias_7 <= 8'h00;
      bias_8 <= 8'h00;
      bias_9 <= 8'h00;
      bias_10 <= 8'h00;
      bias_11 <= 8'h00;
      bias_12 <= 8'h00;
      bias_13 <= 8'h00;
      bias_14 <= 8'h00;
      bias_15 <= 8'h00;
      bias_16 <= 8'h00;
      bias_17 <= 8'h00;
      bias_18 <= 8'h00;
      bias_19 <= 8'h00;
      bias_20 <= 8'h00;
      bias_21 <= 8'h00;
      bias_22 <= 8'h00;
      bias_23 <= 8'h00;
      bias_24 <= 8'h00;
      bias_25 <= 8'h00;
      bias_26 <= 8'h00;
      bias_27 <= 8'h00;
      bias_28 <= 8'h00;
      bias_29 <= 8'h00;
      bias_30 <= 8'h00;
      bias_31 <= 8'h00;
      io_weight_1_delay_1 <= 8'h00;
      io_weight_2_delay_1 <= 8'h00;
      io_weight_2_delay_2 <= 8'h00;
      io_weight_3_delay_1 <= 8'h00;
      io_weight_3_delay_2 <= 8'h00;
      io_weight_3_delay_3 <= 8'h00;
      io_weight_4_delay_1 <= 8'h00;
      io_weight_4_delay_2 <= 8'h00;
      io_weight_4_delay_3 <= 8'h00;
      io_weight_4_delay_4 <= 8'h00;
      io_weight_5_delay_1 <= 8'h00;
      io_weight_5_delay_2 <= 8'h00;
      io_weight_5_delay_3 <= 8'h00;
      io_weight_5_delay_4 <= 8'h00;
      io_weight_5_delay_5 <= 8'h00;
      io_weight_6_delay_1 <= 8'h00;
      io_weight_6_delay_2 <= 8'h00;
      io_weight_6_delay_3 <= 8'h00;
      io_weight_6_delay_4 <= 8'h00;
      io_weight_6_delay_5 <= 8'h00;
      io_weight_6_delay_6 <= 8'h00;
      io_weight_7_delay_1 <= 8'h00;
      io_weight_7_delay_2 <= 8'h00;
      io_weight_7_delay_3 <= 8'h00;
      io_weight_7_delay_4 <= 8'h00;
      io_weight_7_delay_5 <= 8'h00;
      io_weight_7_delay_6 <= 8'h00;
      io_weight_7_delay_7 <= 8'h00;
      io_weight_8_delay_1 <= 8'h00;
      io_weight_8_delay_2 <= 8'h00;
      io_weight_8_delay_3 <= 8'h00;
      io_weight_8_delay_4 <= 8'h00;
      io_weight_8_delay_5 <= 8'h00;
      io_weight_8_delay_6 <= 8'h00;
      io_weight_8_delay_7 <= 8'h00;
      io_weight_8_delay_8 <= 8'h00;
      io_weight_9_delay_1 <= 8'h00;
      io_weight_9_delay_2 <= 8'h00;
      io_weight_9_delay_3 <= 8'h00;
      io_weight_9_delay_4 <= 8'h00;
      io_weight_9_delay_5 <= 8'h00;
      io_weight_9_delay_6 <= 8'h00;
      io_weight_9_delay_7 <= 8'h00;
      io_weight_9_delay_8 <= 8'h00;
      io_weight_9_delay_9 <= 8'h00;
      io_weight_10_delay_1 <= 8'h00;
      io_weight_10_delay_2 <= 8'h00;
      io_weight_10_delay_3 <= 8'h00;
      io_weight_10_delay_4 <= 8'h00;
      io_weight_10_delay_5 <= 8'h00;
      io_weight_10_delay_6 <= 8'h00;
      io_weight_10_delay_7 <= 8'h00;
      io_weight_10_delay_8 <= 8'h00;
      io_weight_10_delay_9 <= 8'h00;
      io_weight_10_delay_10 <= 8'h00;
      io_weight_11_delay_1 <= 8'h00;
      io_weight_11_delay_2 <= 8'h00;
      io_weight_11_delay_3 <= 8'h00;
      io_weight_11_delay_4 <= 8'h00;
      io_weight_11_delay_5 <= 8'h00;
      io_weight_11_delay_6 <= 8'h00;
      io_weight_11_delay_7 <= 8'h00;
      io_weight_11_delay_8 <= 8'h00;
      io_weight_11_delay_9 <= 8'h00;
      io_weight_11_delay_10 <= 8'h00;
      io_weight_11_delay_11 <= 8'h00;
      io_weight_12_delay_1 <= 8'h00;
      io_weight_12_delay_2 <= 8'h00;
      io_weight_12_delay_3 <= 8'h00;
      io_weight_12_delay_4 <= 8'h00;
      io_weight_12_delay_5 <= 8'h00;
      io_weight_12_delay_6 <= 8'h00;
      io_weight_12_delay_7 <= 8'h00;
      io_weight_12_delay_8 <= 8'h00;
      io_weight_12_delay_9 <= 8'h00;
      io_weight_12_delay_10 <= 8'h00;
      io_weight_12_delay_11 <= 8'h00;
      io_weight_12_delay_12 <= 8'h00;
      io_weight_13_delay_1 <= 8'h00;
      io_weight_13_delay_2 <= 8'h00;
      io_weight_13_delay_3 <= 8'h00;
      io_weight_13_delay_4 <= 8'h00;
      io_weight_13_delay_5 <= 8'h00;
      io_weight_13_delay_6 <= 8'h00;
      io_weight_13_delay_7 <= 8'h00;
      io_weight_13_delay_8 <= 8'h00;
      io_weight_13_delay_9 <= 8'h00;
      io_weight_13_delay_10 <= 8'h00;
      io_weight_13_delay_11 <= 8'h00;
      io_weight_13_delay_12 <= 8'h00;
      io_weight_13_delay_13 <= 8'h00;
      io_weight_14_delay_1 <= 8'h00;
      io_weight_14_delay_2 <= 8'h00;
      io_weight_14_delay_3 <= 8'h00;
      io_weight_14_delay_4 <= 8'h00;
      io_weight_14_delay_5 <= 8'h00;
      io_weight_14_delay_6 <= 8'h00;
      io_weight_14_delay_7 <= 8'h00;
      io_weight_14_delay_8 <= 8'h00;
      io_weight_14_delay_9 <= 8'h00;
      io_weight_14_delay_10 <= 8'h00;
      io_weight_14_delay_11 <= 8'h00;
      io_weight_14_delay_12 <= 8'h00;
      io_weight_14_delay_13 <= 8'h00;
      io_weight_14_delay_14 <= 8'h00;
      io_weight_15_delay_1 <= 8'h00;
      io_weight_15_delay_2 <= 8'h00;
      io_weight_15_delay_3 <= 8'h00;
      io_weight_15_delay_4 <= 8'h00;
      io_weight_15_delay_5 <= 8'h00;
      io_weight_15_delay_6 <= 8'h00;
      io_weight_15_delay_7 <= 8'h00;
      io_weight_15_delay_8 <= 8'h00;
      io_weight_15_delay_9 <= 8'h00;
      io_weight_15_delay_10 <= 8'h00;
      io_weight_15_delay_11 <= 8'h00;
      io_weight_15_delay_12 <= 8'h00;
      io_weight_15_delay_13 <= 8'h00;
      io_weight_15_delay_14 <= 8'h00;
      io_weight_15_delay_15 <= 8'h00;
      io_weight_16_delay_1 <= 8'h00;
      io_weight_16_delay_2 <= 8'h00;
      io_weight_16_delay_3 <= 8'h00;
      io_weight_16_delay_4 <= 8'h00;
      io_weight_16_delay_5 <= 8'h00;
      io_weight_16_delay_6 <= 8'h00;
      io_weight_16_delay_7 <= 8'h00;
      io_weight_16_delay_8 <= 8'h00;
      io_weight_16_delay_9 <= 8'h00;
      io_weight_16_delay_10 <= 8'h00;
      io_weight_16_delay_11 <= 8'h00;
      io_weight_16_delay_12 <= 8'h00;
      io_weight_16_delay_13 <= 8'h00;
      io_weight_16_delay_14 <= 8'h00;
      io_weight_16_delay_15 <= 8'h00;
      io_weight_16_delay_16 <= 8'h00;
      io_weight_17_delay_1 <= 8'h00;
      io_weight_17_delay_2 <= 8'h00;
      io_weight_17_delay_3 <= 8'h00;
      io_weight_17_delay_4 <= 8'h00;
      io_weight_17_delay_5 <= 8'h00;
      io_weight_17_delay_6 <= 8'h00;
      io_weight_17_delay_7 <= 8'h00;
      io_weight_17_delay_8 <= 8'h00;
      io_weight_17_delay_9 <= 8'h00;
      io_weight_17_delay_10 <= 8'h00;
      io_weight_17_delay_11 <= 8'h00;
      io_weight_17_delay_12 <= 8'h00;
      io_weight_17_delay_13 <= 8'h00;
      io_weight_17_delay_14 <= 8'h00;
      io_weight_17_delay_15 <= 8'h00;
      io_weight_17_delay_16 <= 8'h00;
      io_weight_17_delay_17 <= 8'h00;
      io_weight_18_delay_1 <= 8'h00;
      io_weight_18_delay_2 <= 8'h00;
      io_weight_18_delay_3 <= 8'h00;
      io_weight_18_delay_4 <= 8'h00;
      io_weight_18_delay_5 <= 8'h00;
      io_weight_18_delay_6 <= 8'h00;
      io_weight_18_delay_7 <= 8'h00;
      io_weight_18_delay_8 <= 8'h00;
      io_weight_18_delay_9 <= 8'h00;
      io_weight_18_delay_10 <= 8'h00;
      io_weight_18_delay_11 <= 8'h00;
      io_weight_18_delay_12 <= 8'h00;
      io_weight_18_delay_13 <= 8'h00;
      io_weight_18_delay_14 <= 8'h00;
      io_weight_18_delay_15 <= 8'h00;
      io_weight_18_delay_16 <= 8'h00;
      io_weight_18_delay_17 <= 8'h00;
      io_weight_18_delay_18 <= 8'h00;
      io_weight_19_delay_1 <= 8'h00;
      io_weight_19_delay_2 <= 8'h00;
      io_weight_19_delay_3 <= 8'h00;
      io_weight_19_delay_4 <= 8'h00;
      io_weight_19_delay_5 <= 8'h00;
      io_weight_19_delay_6 <= 8'h00;
      io_weight_19_delay_7 <= 8'h00;
      io_weight_19_delay_8 <= 8'h00;
      io_weight_19_delay_9 <= 8'h00;
      io_weight_19_delay_10 <= 8'h00;
      io_weight_19_delay_11 <= 8'h00;
      io_weight_19_delay_12 <= 8'h00;
      io_weight_19_delay_13 <= 8'h00;
      io_weight_19_delay_14 <= 8'h00;
      io_weight_19_delay_15 <= 8'h00;
      io_weight_19_delay_16 <= 8'h00;
      io_weight_19_delay_17 <= 8'h00;
      io_weight_19_delay_18 <= 8'h00;
      io_weight_19_delay_19 <= 8'h00;
      io_weight_20_delay_1 <= 8'h00;
      io_weight_20_delay_2 <= 8'h00;
      io_weight_20_delay_3 <= 8'h00;
      io_weight_20_delay_4 <= 8'h00;
      io_weight_20_delay_5 <= 8'h00;
      io_weight_20_delay_6 <= 8'h00;
      io_weight_20_delay_7 <= 8'h00;
      io_weight_20_delay_8 <= 8'h00;
      io_weight_20_delay_9 <= 8'h00;
      io_weight_20_delay_10 <= 8'h00;
      io_weight_20_delay_11 <= 8'h00;
      io_weight_20_delay_12 <= 8'h00;
      io_weight_20_delay_13 <= 8'h00;
      io_weight_20_delay_14 <= 8'h00;
      io_weight_20_delay_15 <= 8'h00;
      io_weight_20_delay_16 <= 8'h00;
      io_weight_20_delay_17 <= 8'h00;
      io_weight_20_delay_18 <= 8'h00;
      io_weight_20_delay_19 <= 8'h00;
      io_weight_20_delay_20 <= 8'h00;
      io_weight_21_delay_1 <= 8'h00;
      io_weight_21_delay_2 <= 8'h00;
      io_weight_21_delay_3 <= 8'h00;
      io_weight_21_delay_4 <= 8'h00;
      io_weight_21_delay_5 <= 8'h00;
      io_weight_21_delay_6 <= 8'h00;
      io_weight_21_delay_7 <= 8'h00;
      io_weight_21_delay_8 <= 8'h00;
      io_weight_21_delay_9 <= 8'h00;
      io_weight_21_delay_10 <= 8'h00;
      io_weight_21_delay_11 <= 8'h00;
      io_weight_21_delay_12 <= 8'h00;
      io_weight_21_delay_13 <= 8'h00;
      io_weight_21_delay_14 <= 8'h00;
      io_weight_21_delay_15 <= 8'h00;
      io_weight_21_delay_16 <= 8'h00;
      io_weight_21_delay_17 <= 8'h00;
      io_weight_21_delay_18 <= 8'h00;
      io_weight_21_delay_19 <= 8'h00;
      io_weight_21_delay_20 <= 8'h00;
      io_weight_21_delay_21 <= 8'h00;
      io_weight_22_delay_1 <= 8'h00;
      io_weight_22_delay_2 <= 8'h00;
      io_weight_22_delay_3 <= 8'h00;
      io_weight_22_delay_4 <= 8'h00;
      io_weight_22_delay_5 <= 8'h00;
      io_weight_22_delay_6 <= 8'h00;
      io_weight_22_delay_7 <= 8'h00;
      io_weight_22_delay_8 <= 8'h00;
      io_weight_22_delay_9 <= 8'h00;
      io_weight_22_delay_10 <= 8'h00;
      io_weight_22_delay_11 <= 8'h00;
      io_weight_22_delay_12 <= 8'h00;
      io_weight_22_delay_13 <= 8'h00;
      io_weight_22_delay_14 <= 8'h00;
      io_weight_22_delay_15 <= 8'h00;
      io_weight_22_delay_16 <= 8'h00;
      io_weight_22_delay_17 <= 8'h00;
      io_weight_22_delay_18 <= 8'h00;
      io_weight_22_delay_19 <= 8'h00;
      io_weight_22_delay_20 <= 8'h00;
      io_weight_22_delay_21 <= 8'h00;
      io_weight_22_delay_22 <= 8'h00;
      io_weight_23_delay_1 <= 8'h00;
      io_weight_23_delay_2 <= 8'h00;
      io_weight_23_delay_3 <= 8'h00;
      io_weight_23_delay_4 <= 8'h00;
      io_weight_23_delay_5 <= 8'h00;
      io_weight_23_delay_6 <= 8'h00;
      io_weight_23_delay_7 <= 8'h00;
      io_weight_23_delay_8 <= 8'h00;
      io_weight_23_delay_9 <= 8'h00;
      io_weight_23_delay_10 <= 8'h00;
      io_weight_23_delay_11 <= 8'h00;
      io_weight_23_delay_12 <= 8'h00;
      io_weight_23_delay_13 <= 8'h00;
      io_weight_23_delay_14 <= 8'h00;
      io_weight_23_delay_15 <= 8'h00;
      io_weight_23_delay_16 <= 8'h00;
      io_weight_23_delay_17 <= 8'h00;
      io_weight_23_delay_18 <= 8'h00;
      io_weight_23_delay_19 <= 8'h00;
      io_weight_23_delay_20 <= 8'h00;
      io_weight_23_delay_21 <= 8'h00;
      io_weight_23_delay_22 <= 8'h00;
      io_weight_23_delay_23 <= 8'h00;
      io_weight_24_delay_1 <= 8'h00;
      io_weight_24_delay_2 <= 8'h00;
      io_weight_24_delay_3 <= 8'h00;
      io_weight_24_delay_4 <= 8'h00;
      io_weight_24_delay_5 <= 8'h00;
      io_weight_24_delay_6 <= 8'h00;
      io_weight_24_delay_7 <= 8'h00;
      io_weight_24_delay_8 <= 8'h00;
      io_weight_24_delay_9 <= 8'h00;
      io_weight_24_delay_10 <= 8'h00;
      io_weight_24_delay_11 <= 8'h00;
      io_weight_24_delay_12 <= 8'h00;
      io_weight_24_delay_13 <= 8'h00;
      io_weight_24_delay_14 <= 8'h00;
      io_weight_24_delay_15 <= 8'h00;
      io_weight_24_delay_16 <= 8'h00;
      io_weight_24_delay_17 <= 8'h00;
      io_weight_24_delay_18 <= 8'h00;
      io_weight_24_delay_19 <= 8'h00;
      io_weight_24_delay_20 <= 8'h00;
      io_weight_24_delay_21 <= 8'h00;
      io_weight_24_delay_22 <= 8'h00;
      io_weight_24_delay_23 <= 8'h00;
      io_weight_24_delay_24 <= 8'h00;
      io_weight_25_delay_1 <= 8'h00;
      io_weight_25_delay_2 <= 8'h00;
      io_weight_25_delay_3 <= 8'h00;
      io_weight_25_delay_4 <= 8'h00;
      io_weight_25_delay_5 <= 8'h00;
      io_weight_25_delay_6 <= 8'h00;
      io_weight_25_delay_7 <= 8'h00;
      io_weight_25_delay_8 <= 8'h00;
      io_weight_25_delay_9 <= 8'h00;
      io_weight_25_delay_10 <= 8'h00;
      io_weight_25_delay_11 <= 8'h00;
      io_weight_25_delay_12 <= 8'h00;
      io_weight_25_delay_13 <= 8'h00;
      io_weight_25_delay_14 <= 8'h00;
      io_weight_25_delay_15 <= 8'h00;
      io_weight_25_delay_16 <= 8'h00;
      io_weight_25_delay_17 <= 8'h00;
      io_weight_25_delay_18 <= 8'h00;
      io_weight_25_delay_19 <= 8'h00;
      io_weight_25_delay_20 <= 8'h00;
      io_weight_25_delay_21 <= 8'h00;
      io_weight_25_delay_22 <= 8'h00;
      io_weight_25_delay_23 <= 8'h00;
      io_weight_25_delay_24 <= 8'h00;
      io_weight_25_delay_25 <= 8'h00;
      io_weight_26_delay_1 <= 8'h00;
      io_weight_26_delay_2 <= 8'h00;
      io_weight_26_delay_3 <= 8'h00;
      io_weight_26_delay_4 <= 8'h00;
      io_weight_26_delay_5 <= 8'h00;
      io_weight_26_delay_6 <= 8'h00;
      io_weight_26_delay_7 <= 8'h00;
      io_weight_26_delay_8 <= 8'h00;
      io_weight_26_delay_9 <= 8'h00;
      io_weight_26_delay_10 <= 8'h00;
      io_weight_26_delay_11 <= 8'h00;
      io_weight_26_delay_12 <= 8'h00;
      io_weight_26_delay_13 <= 8'h00;
      io_weight_26_delay_14 <= 8'h00;
      io_weight_26_delay_15 <= 8'h00;
      io_weight_26_delay_16 <= 8'h00;
      io_weight_26_delay_17 <= 8'h00;
      io_weight_26_delay_18 <= 8'h00;
      io_weight_26_delay_19 <= 8'h00;
      io_weight_26_delay_20 <= 8'h00;
      io_weight_26_delay_21 <= 8'h00;
      io_weight_26_delay_22 <= 8'h00;
      io_weight_26_delay_23 <= 8'h00;
      io_weight_26_delay_24 <= 8'h00;
      io_weight_26_delay_25 <= 8'h00;
      io_weight_26_delay_26 <= 8'h00;
      io_weight_27_delay_1 <= 8'h00;
      io_weight_27_delay_2 <= 8'h00;
      io_weight_27_delay_3 <= 8'h00;
      io_weight_27_delay_4 <= 8'h00;
      io_weight_27_delay_5 <= 8'h00;
      io_weight_27_delay_6 <= 8'h00;
      io_weight_27_delay_7 <= 8'h00;
      io_weight_27_delay_8 <= 8'h00;
      io_weight_27_delay_9 <= 8'h00;
      io_weight_27_delay_10 <= 8'h00;
      io_weight_27_delay_11 <= 8'h00;
      io_weight_27_delay_12 <= 8'h00;
      io_weight_27_delay_13 <= 8'h00;
      io_weight_27_delay_14 <= 8'h00;
      io_weight_27_delay_15 <= 8'h00;
      io_weight_27_delay_16 <= 8'h00;
      io_weight_27_delay_17 <= 8'h00;
      io_weight_27_delay_18 <= 8'h00;
      io_weight_27_delay_19 <= 8'h00;
      io_weight_27_delay_20 <= 8'h00;
      io_weight_27_delay_21 <= 8'h00;
      io_weight_27_delay_22 <= 8'h00;
      io_weight_27_delay_23 <= 8'h00;
      io_weight_27_delay_24 <= 8'h00;
      io_weight_27_delay_25 <= 8'h00;
      io_weight_27_delay_26 <= 8'h00;
      io_weight_27_delay_27 <= 8'h00;
      io_weight_28_delay_1 <= 8'h00;
      io_weight_28_delay_2 <= 8'h00;
      io_weight_28_delay_3 <= 8'h00;
      io_weight_28_delay_4 <= 8'h00;
      io_weight_28_delay_5 <= 8'h00;
      io_weight_28_delay_6 <= 8'h00;
      io_weight_28_delay_7 <= 8'h00;
      io_weight_28_delay_8 <= 8'h00;
      io_weight_28_delay_9 <= 8'h00;
      io_weight_28_delay_10 <= 8'h00;
      io_weight_28_delay_11 <= 8'h00;
      io_weight_28_delay_12 <= 8'h00;
      io_weight_28_delay_13 <= 8'h00;
      io_weight_28_delay_14 <= 8'h00;
      io_weight_28_delay_15 <= 8'h00;
      io_weight_28_delay_16 <= 8'h00;
      io_weight_28_delay_17 <= 8'h00;
      io_weight_28_delay_18 <= 8'h00;
      io_weight_28_delay_19 <= 8'h00;
      io_weight_28_delay_20 <= 8'h00;
      io_weight_28_delay_21 <= 8'h00;
      io_weight_28_delay_22 <= 8'h00;
      io_weight_28_delay_23 <= 8'h00;
      io_weight_28_delay_24 <= 8'h00;
      io_weight_28_delay_25 <= 8'h00;
      io_weight_28_delay_26 <= 8'h00;
      io_weight_28_delay_27 <= 8'h00;
      io_weight_28_delay_28 <= 8'h00;
      io_weight_29_delay_1 <= 8'h00;
      io_weight_29_delay_2 <= 8'h00;
      io_weight_29_delay_3 <= 8'h00;
      io_weight_29_delay_4 <= 8'h00;
      io_weight_29_delay_5 <= 8'h00;
      io_weight_29_delay_6 <= 8'h00;
      io_weight_29_delay_7 <= 8'h00;
      io_weight_29_delay_8 <= 8'h00;
      io_weight_29_delay_9 <= 8'h00;
      io_weight_29_delay_10 <= 8'h00;
      io_weight_29_delay_11 <= 8'h00;
      io_weight_29_delay_12 <= 8'h00;
      io_weight_29_delay_13 <= 8'h00;
      io_weight_29_delay_14 <= 8'h00;
      io_weight_29_delay_15 <= 8'h00;
      io_weight_29_delay_16 <= 8'h00;
      io_weight_29_delay_17 <= 8'h00;
      io_weight_29_delay_18 <= 8'h00;
      io_weight_29_delay_19 <= 8'h00;
      io_weight_29_delay_20 <= 8'h00;
      io_weight_29_delay_21 <= 8'h00;
      io_weight_29_delay_22 <= 8'h00;
      io_weight_29_delay_23 <= 8'h00;
      io_weight_29_delay_24 <= 8'h00;
      io_weight_29_delay_25 <= 8'h00;
      io_weight_29_delay_26 <= 8'h00;
      io_weight_29_delay_27 <= 8'h00;
      io_weight_29_delay_28 <= 8'h00;
      io_weight_29_delay_29 <= 8'h00;
      io_weight_30_delay_1 <= 8'h00;
      io_weight_30_delay_2 <= 8'h00;
      io_weight_30_delay_3 <= 8'h00;
      io_weight_30_delay_4 <= 8'h00;
      io_weight_30_delay_5 <= 8'h00;
      io_weight_30_delay_6 <= 8'h00;
      io_weight_30_delay_7 <= 8'h00;
      io_weight_30_delay_8 <= 8'h00;
      io_weight_30_delay_9 <= 8'h00;
      io_weight_30_delay_10 <= 8'h00;
      io_weight_30_delay_11 <= 8'h00;
      io_weight_30_delay_12 <= 8'h00;
      io_weight_30_delay_13 <= 8'h00;
      io_weight_30_delay_14 <= 8'h00;
      io_weight_30_delay_15 <= 8'h00;
      io_weight_30_delay_16 <= 8'h00;
      io_weight_30_delay_17 <= 8'h00;
      io_weight_30_delay_18 <= 8'h00;
      io_weight_30_delay_19 <= 8'h00;
      io_weight_30_delay_20 <= 8'h00;
      io_weight_30_delay_21 <= 8'h00;
      io_weight_30_delay_22 <= 8'h00;
      io_weight_30_delay_23 <= 8'h00;
      io_weight_30_delay_24 <= 8'h00;
      io_weight_30_delay_25 <= 8'h00;
      io_weight_30_delay_26 <= 8'h00;
      io_weight_30_delay_27 <= 8'h00;
      io_weight_30_delay_28 <= 8'h00;
      io_weight_30_delay_29 <= 8'h00;
      io_weight_30_delay_30 <= 8'h00;
      io_weight_31_delay_1 <= 8'h00;
      io_weight_31_delay_2 <= 8'h00;
      io_weight_31_delay_3 <= 8'h00;
      io_weight_31_delay_4 <= 8'h00;
      io_weight_31_delay_5 <= 8'h00;
      io_weight_31_delay_6 <= 8'h00;
      io_weight_31_delay_7 <= 8'h00;
      io_weight_31_delay_8 <= 8'h00;
      io_weight_31_delay_9 <= 8'h00;
      io_weight_31_delay_10 <= 8'h00;
      io_weight_31_delay_11 <= 8'h00;
      io_weight_31_delay_12 <= 8'h00;
      io_weight_31_delay_13 <= 8'h00;
      io_weight_31_delay_14 <= 8'h00;
      io_weight_31_delay_15 <= 8'h00;
      io_weight_31_delay_16 <= 8'h00;
      io_weight_31_delay_17 <= 8'h00;
      io_weight_31_delay_18 <= 8'h00;
      io_weight_31_delay_19 <= 8'h00;
      io_weight_31_delay_20 <= 8'h00;
      io_weight_31_delay_21 <= 8'h00;
      io_weight_31_delay_22 <= 8'h00;
      io_weight_31_delay_23 <= 8'h00;
      io_weight_31_delay_24 <= 8'h00;
      io_weight_31_delay_25 <= 8'h00;
      io_weight_31_delay_26 <= 8'h00;
      io_weight_31_delay_27 <= 8'h00;
      io_weight_31_delay_28 <= 8'h00;
      io_weight_31_delay_29 <= 8'h00;
      io_weight_31_delay_30 <= 8'h00;
      io_weight_31_delay_31 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_9 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_10 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_11 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_12 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_13 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_14 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_15 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_16 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_17 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_18 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_19 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_20 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_21 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_22 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_23 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_24 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_25 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_26 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_27 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_28 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_29 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_30 <= 8'h00;
      toplevel_mac_0_31_io_macOut_delay_31 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_9 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_10 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_11 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_12 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_13 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_14 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_15 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_16 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_17 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_18 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_19 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_20 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_21 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_22 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_23 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_24 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_25 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_26 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_27 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_28 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_29 <= 8'h00;
      toplevel_mac_1_31_io_macOut_delay_30 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_9 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_10 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_11 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_12 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_13 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_14 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_15 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_16 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_17 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_18 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_19 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_20 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_21 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_22 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_23 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_24 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_25 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_26 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_27 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_28 <= 8'h00;
      toplevel_mac_2_31_io_macOut_delay_29 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_9 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_10 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_11 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_12 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_13 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_14 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_15 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_16 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_17 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_18 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_19 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_20 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_21 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_22 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_23 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_24 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_25 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_26 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_27 <= 8'h00;
      toplevel_mac_3_31_io_macOut_delay_28 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_9 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_10 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_11 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_12 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_13 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_14 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_15 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_16 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_17 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_18 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_19 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_20 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_21 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_22 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_23 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_24 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_25 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_26 <= 8'h00;
      toplevel_mac_4_31_io_macOut_delay_27 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_9 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_10 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_11 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_12 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_13 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_14 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_15 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_16 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_17 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_18 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_19 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_20 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_21 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_22 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_23 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_24 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_25 <= 8'h00;
      toplevel_mac_5_31_io_macOut_delay_26 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_9 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_10 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_11 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_12 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_13 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_14 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_15 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_16 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_17 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_18 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_19 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_20 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_21 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_22 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_23 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_24 <= 8'h00;
      toplevel_mac_6_31_io_macOut_delay_25 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_9 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_10 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_11 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_12 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_13 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_14 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_15 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_16 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_17 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_18 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_19 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_20 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_21 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_22 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_23 <= 8'h00;
      toplevel_mac_7_31_io_macOut_delay_24 <= 8'h00;
      toplevel_mac_8_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_8_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_8_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_8_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_8_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_8_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_8_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_8_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_8_31_io_macOut_delay_9 <= 8'h00;
      toplevel_mac_8_31_io_macOut_delay_10 <= 8'h00;
      toplevel_mac_8_31_io_macOut_delay_11 <= 8'h00;
      toplevel_mac_8_31_io_macOut_delay_12 <= 8'h00;
      toplevel_mac_8_31_io_macOut_delay_13 <= 8'h00;
      toplevel_mac_8_31_io_macOut_delay_14 <= 8'h00;
      toplevel_mac_8_31_io_macOut_delay_15 <= 8'h00;
      toplevel_mac_8_31_io_macOut_delay_16 <= 8'h00;
      toplevel_mac_8_31_io_macOut_delay_17 <= 8'h00;
      toplevel_mac_8_31_io_macOut_delay_18 <= 8'h00;
      toplevel_mac_8_31_io_macOut_delay_19 <= 8'h00;
      toplevel_mac_8_31_io_macOut_delay_20 <= 8'h00;
      toplevel_mac_8_31_io_macOut_delay_21 <= 8'h00;
      toplevel_mac_8_31_io_macOut_delay_22 <= 8'h00;
      toplevel_mac_8_31_io_macOut_delay_23 <= 8'h00;
      toplevel_mac_9_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_9_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_9_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_9_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_9_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_9_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_9_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_9_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_9_31_io_macOut_delay_9 <= 8'h00;
      toplevel_mac_9_31_io_macOut_delay_10 <= 8'h00;
      toplevel_mac_9_31_io_macOut_delay_11 <= 8'h00;
      toplevel_mac_9_31_io_macOut_delay_12 <= 8'h00;
      toplevel_mac_9_31_io_macOut_delay_13 <= 8'h00;
      toplevel_mac_9_31_io_macOut_delay_14 <= 8'h00;
      toplevel_mac_9_31_io_macOut_delay_15 <= 8'h00;
      toplevel_mac_9_31_io_macOut_delay_16 <= 8'h00;
      toplevel_mac_9_31_io_macOut_delay_17 <= 8'h00;
      toplevel_mac_9_31_io_macOut_delay_18 <= 8'h00;
      toplevel_mac_9_31_io_macOut_delay_19 <= 8'h00;
      toplevel_mac_9_31_io_macOut_delay_20 <= 8'h00;
      toplevel_mac_9_31_io_macOut_delay_21 <= 8'h00;
      toplevel_mac_9_31_io_macOut_delay_22 <= 8'h00;
      toplevel_mac_10_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_10_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_10_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_10_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_10_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_10_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_10_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_10_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_10_31_io_macOut_delay_9 <= 8'h00;
      toplevel_mac_10_31_io_macOut_delay_10 <= 8'h00;
      toplevel_mac_10_31_io_macOut_delay_11 <= 8'h00;
      toplevel_mac_10_31_io_macOut_delay_12 <= 8'h00;
      toplevel_mac_10_31_io_macOut_delay_13 <= 8'h00;
      toplevel_mac_10_31_io_macOut_delay_14 <= 8'h00;
      toplevel_mac_10_31_io_macOut_delay_15 <= 8'h00;
      toplevel_mac_10_31_io_macOut_delay_16 <= 8'h00;
      toplevel_mac_10_31_io_macOut_delay_17 <= 8'h00;
      toplevel_mac_10_31_io_macOut_delay_18 <= 8'h00;
      toplevel_mac_10_31_io_macOut_delay_19 <= 8'h00;
      toplevel_mac_10_31_io_macOut_delay_20 <= 8'h00;
      toplevel_mac_10_31_io_macOut_delay_21 <= 8'h00;
      toplevel_mac_11_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_11_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_11_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_11_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_11_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_11_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_11_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_11_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_11_31_io_macOut_delay_9 <= 8'h00;
      toplevel_mac_11_31_io_macOut_delay_10 <= 8'h00;
      toplevel_mac_11_31_io_macOut_delay_11 <= 8'h00;
      toplevel_mac_11_31_io_macOut_delay_12 <= 8'h00;
      toplevel_mac_11_31_io_macOut_delay_13 <= 8'h00;
      toplevel_mac_11_31_io_macOut_delay_14 <= 8'h00;
      toplevel_mac_11_31_io_macOut_delay_15 <= 8'h00;
      toplevel_mac_11_31_io_macOut_delay_16 <= 8'h00;
      toplevel_mac_11_31_io_macOut_delay_17 <= 8'h00;
      toplevel_mac_11_31_io_macOut_delay_18 <= 8'h00;
      toplevel_mac_11_31_io_macOut_delay_19 <= 8'h00;
      toplevel_mac_11_31_io_macOut_delay_20 <= 8'h00;
      toplevel_mac_12_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_12_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_12_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_12_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_12_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_12_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_12_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_12_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_12_31_io_macOut_delay_9 <= 8'h00;
      toplevel_mac_12_31_io_macOut_delay_10 <= 8'h00;
      toplevel_mac_12_31_io_macOut_delay_11 <= 8'h00;
      toplevel_mac_12_31_io_macOut_delay_12 <= 8'h00;
      toplevel_mac_12_31_io_macOut_delay_13 <= 8'h00;
      toplevel_mac_12_31_io_macOut_delay_14 <= 8'h00;
      toplevel_mac_12_31_io_macOut_delay_15 <= 8'h00;
      toplevel_mac_12_31_io_macOut_delay_16 <= 8'h00;
      toplevel_mac_12_31_io_macOut_delay_17 <= 8'h00;
      toplevel_mac_12_31_io_macOut_delay_18 <= 8'h00;
      toplevel_mac_12_31_io_macOut_delay_19 <= 8'h00;
      toplevel_mac_13_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_13_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_13_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_13_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_13_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_13_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_13_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_13_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_13_31_io_macOut_delay_9 <= 8'h00;
      toplevel_mac_13_31_io_macOut_delay_10 <= 8'h00;
      toplevel_mac_13_31_io_macOut_delay_11 <= 8'h00;
      toplevel_mac_13_31_io_macOut_delay_12 <= 8'h00;
      toplevel_mac_13_31_io_macOut_delay_13 <= 8'h00;
      toplevel_mac_13_31_io_macOut_delay_14 <= 8'h00;
      toplevel_mac_13_31_io_macOut_delay_15 <= 8'h00;
      toplevel_mac_13_31_io_macOut_delay_16 <= 8'h00;
      toplevel_mac_13_31_io_macOut_delay_17 <= 8'h00;
      toplevel_mac_13_31_io_macOut_delay_18 <= 8'h00;
      toplevel_mac_14_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_14_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_14_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_14_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_14_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_14_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_14_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_14_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_14_31_io_macOut_delay_9 <= 8'h00;
      toplevel_mac_14_31_io_macOut_delay_10 <= 8'h00;
      toplevel_mac_14_31_io_macOut_delay_11 <= 8'h00;
      toplevel_mac_14_31_io_macOut_delay_12 <= 8'h00;
      toplevel_mac_14_31_io_macOut_delay_13 <= 8'h00;
      toplevel_mac_14_31_io_macOut_delay_14 <= 8'h00;
      toplevel_mac_14_31_io_macOut_delay_15 <= 8'h00;
      toplevel_mac_14_31_io_macOut_delay_16 <= 8'h00;
      toplevel_mac_14_31_io_macOut_delay_17 <= 8'h00;
      toplevel_mac_15_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_15_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_15_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_15_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_15_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_15_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_15_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_15_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_15_31_io_macOut_delay_9 <= 8'h00;
      toplevel_mac_15_31_io_macOut_delay_10 <= 8'h00;
      toplevel_mac_15_31_io_macOut_delay_11 <= 8'h00;
      toplevel_mac_15_31_io_macOut_delay_12 <= 8'h00;
      toplevel_mac_15_31_io_macOut_delay_13 <= 8'h00;
      toplevel_mac_15_31_io_macOut_delay_14 <= 8'h00;
      toplevel_mac_15_31_io_macOut_delay_15 <= 8'h00;
      toplevel_mac_15_31_io_macOut_delay_16 <= 8'h00;
      toplevel_mac_16_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_16_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_16_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_16_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_16_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_16_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_16_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_16_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_16_31_io_macOut_delay_9 <= 8'h00;
      toplevel_mac_16_31_io_macOut_delay_10 <= 8'h00;
      toplevel_mac_16_31_io_macOut_delay_11 <= 8'h00;
      toplevel_mac_16_31_io_macOut_delay_12 <= 8'h00;
      toplevel_mac_16_31_io_macOut_delay_13 <= 8'h00;
      toplevel_mac_16_31_io_macOut_delay_14 <= 8'h00;
      toplevel_mac_16_31_io_macOut_delay_15 <= 8'h00;
      toplevel_mac_17_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_17_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_17_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_17_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_17_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_17_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_17_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_17_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_17_31_io_macOut_delay_9 <= 8'h00;
      toplevel_mac_17_31_io_macOut_delay_10 <= 8'h00;
      toplevel_mac_17_31_io_macOut_delay_11 <= 8'h00;
      toplevel_mac_17_31_io_macOut_delay_12 <= 8'h00;
      toplevel_mac_17_31_io_macOut_delay_13 <= 8'h00;
      toplevel_mac_17_31_io_macOut_delay_14 <= 8'h00;
      toplevel_mac_18_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_18_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_18_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_18_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_18_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_18_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_18_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_18_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_18_31_io_macOut_delay_9 <= 8'h00;
      toplevel_mac_18_31_io_macOut_delay_10 <= 8'h00;
      toplevel_mac_18_31_io_macOut_delay_11 <= 8'h00;
      toplevel_mac_18_31_io_macOut_delay_12 <= 8'h00;
      toplevel_mac_18_31_io_macOut_delay_13 <= 8'h00;
      toplevel_mac_19_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_19_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_19_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_19_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_19_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_19_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_19_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_19_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_19_31_io_macOut_delay_9 <= 8'h00;
      toplevel_mac_19_31_io_macOut_delay_10 <= 8'h00;
      toplevel_mac_19_31_io_macOut_delay_11 <= 8'h00;
      toplevel_mac_19_31_io_macOut_delay_12 <= 8'h00;
      toplevel_mac_20_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_20_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_20_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_20_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_20_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_20_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_20_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_20_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_20_31_io_macOut_delay_9 <= 8'h00;
      toplevel_mac_20_31_io_macOut_delay_10 <= 8'h00;
      toplevel_mac_20_31_io_macOut_delay_11 <= 8'h00;
      toplevel_mac_21_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_21_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_21_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_21_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_21_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_21_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_21_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_21_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_21_31_io_macOut_delay_9 <= 8'h00;
      toplevel_mac_21_31_io_macOut_delay_10 <= 8'h00;
      toplevel_mac_22_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_22_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_22_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_22_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_22_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_22_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_22_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_22_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_22_31_io_macOut_delay_9 <= 8'h00;
      toplevel_mac_23_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_23_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_23_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_23_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_23_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_23_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_23_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_23_31_io_macOut_delay_8 <= 8'h00;
      toplevel_mac_24_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_24_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_24_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_24_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_24_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_24_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_24_31_io_macOut_delay_7 <= 8'h00;
      toplevel_mac_25_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_25_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_25_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_25_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_25_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_25_31_io_macOut_delay_6 <= 8'h00;
      toplevel_mac_26_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_26_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_26_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_26_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_26_31_io_macOut_delay_5 <= 8'h00;
      toplevel_mac_27_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_27_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_27_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_27_31_io_macOut_delay_4 <= 8'h00;
      toplevel_mac_28_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_28_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_28_31_io_macOut_delay_3 <= 8'h00;
      toplevel_mac_29_31_io_macOut_delay_1 <= 8'h00;
      toplevel_mac_29_31_io_macOut_delay_2 <= 8'h00;
      toplevel_mac_30_31_io_macOut_delay_1 <= 8'h00;
    end else begin
      if(io_load) begin
        bias_0 <= io_activation_0;
        bias_1 <= io_activation_1;
        bias_2 <= io_activation_2;
        bias_3 <= io_activation_3;
        bias_4 <= io_activation_4;
        bias_5 <= io_activation_5;
        bias_6 <= io_activation_6;
        bias_7 <= io_activation_7;
        bias_8 <= io_activation_8;
        bias_9 <= io_activation_9;
        bias_10 <= io_activation_10;
        bias_11 <= io_activation_11;
        bias_12 <= io_activation_12;
        bias_13 <= io_activation_13;
        bias_14 <= io_activation_14;
        bias_15 <= io_activation_15;
        bias_16 <= io_activation_16;
        bias_17 <= io_activation_17;
        bias_18 <= io_activation_18;
        bias_19 <= io_activation_19;
        bias_20 <= io_activation_20;
        bias_21 <= io_activation_21;
        bias_22 <= io_activation_22;
        bias_23 <= io_activation_23;
        bias_24 <= io_activation_24;
        bias_25 <= io_activation_25;
        bias_26 <= io_activation_26;
        bias_27 <= io_activation_27;
        bias_28 <= io_activation_28;
        bias_29 <= io_activation_29;
        bias_30 <= io_activation_30;
        bias_31 <= io_activation_31;
      end
      io_weight_1_delay_1 <= io_weight_1;
      io_weight_2_delay_1 <= io_weight_2;
      io_weight_2_delay_2 <= io_weight_2_delay_1;
      io_weight_3_delay_1 <= io_weight_3;
      io_weight_3_delay_2 <= io_weight_3_delay_1;
      io_weight_3_delay_3 <= io_weight_3_delay_2;
      io_weight_4_delay_1 <= io_weight_4;
      io_weight_4_delay_2 <= io_weight_4_delay_1;
      io_weight_4_delay_3 <= io_weight_4_delay_2;
      io_weight_4_delay_4 <= io_weight_4_delay_3;
      io_weight_5_delay_1 <= io_weight_5;
      io_weight_5_delay_2 <= io_weight_5_delay_1;
      io_weight_5_delay_3 <= io_weight_5_delay_2;
      io_weight_5_delay_4 <= io_weight_5_delay_3;
      io_weight_5_delay_5 <= io_weight_5_delay_4;
      io_weight_6_delay_1 <= io_weight_6;
      io_weight_6_delay_2 <= io_weight_6_delay_1;
      io_weight_6_delay_3 <= io_weight_6_delay_2;
      io_weight_6_delay_4 <= io_weight_6_delay_3;
      io_weight_6_delay_5 <= io_weight_6_delay_4;
      io_weight_6_delay_6 <= io_weight_6_delay_5;
      io_weight_7_delay_1 <= io_weight_7;
      io_weight_7_delay_2 <= io_weight_7_delay_1;
      io_weight_7_delay_3 <= io_weight_7_delay_2;
      io_weight_7_delay_4 <= io_weight_7_delay_3;
      io_weight_7_delay_5 <= io_weight_7_delay_4;
      io_weight_7_delay_6 <= io_weight_7_delay_5;
      io_weight_7_delay_7 <= io_weight_7_delay_6;
      io_weight_8_delay_1 <= io_weight_8;
      io_weight_8_delay_2 <= io_weight_8_delay_1;
      io_weight_8_delay_3 <= io_weight_8_delay_2;
      io_weight_8_delay_4 <= io_weight_8_delay_3;
      io_weight_8_delay_5 <= io_weight_8_delay_4;
      io_weight_8_delay_6 <= io_weight_8_delay_5;
      io_weight_8_delay_7 <= io_weight_8_delay_6;
      io_weight_8_delay_8 <= io_weight_8_delay_7;
      io_weight_9_delay_1 <= io_weight_9;
      io_weight_9_delay_2 <= io_weight_9_delay_1;
      io_weight_9_delay_3 <= io_weight_9_delay_2;
      io_weight_9_delay_4 <= io_weight_9_delay_3;
      io_weight_9_delay_5 <= io_weight_9_delay_4;
      io_weight_9_delay_6 <= io_weight_9_delay_5;
      io_weight_9_delay_7 <= io_weight_9_delay_6;
      io_weight_9_delay_8 <= io_weight_9_delay_7;
      io_weight_9_delay_9 <= io_weight_9_delay_8;
      io_weight_10_delay_1 <= io_weight_10;
      io_weight_10_delay_2 <= io_weight_10_delay_1;
      io_weight_10_delay_3 <= io_weight_10_delay_2;
      io_weight_10_delay_4 <= io_weight_10_delay_3;
      io_weight_10_delay_5 <= io_weight_10_delay_4;
      io_weight_10_delay_6 <= io_weight_10_delay_5;
      io_weight_10_delay_7 <= io_weight_10_delay_6;
      io_weight_10_delay_8 <= io_weight_10_delay_7;
      io_weight_10_delay_9 <= io_weight_10_delay_8;
      io_weight_10_delay_10 <= io_weight_10_delay_9;
      io_weight_11_delay_1 <= io_weight_11;
      io_weight_11_delay_2 <= io_weight_11_delay_1;
      io_weight_11_delay_3 <= io_weight_11_delay_2;
      io_weight_11_delay_4 <= io_weight_11_delay_3;
      io_weight_11_delay_5 <= io_weight_11_delay_4;
      io_weight_11_delay_6 <= io_weight_11_delay_5;
      io_weight_11_delay_7 <= io_weight_11_delay_6;
      io_weight_11_delay_8 <= io_weight_11_delay_7;
      io_weight_11_delay_9 <= io_weight_11_delay_8;
      io_weight_11_delay_10 <= io_weight_11_delay_9;
      io_weight_11_delay_11 <= io_weight_11_delay_10;
      io_weight_12_delay_1 <= io_weight_12;
      io_weight_12_delay_2 <= io_weight_12_delay_1;
      io_weight_12_delay_3 <= io_weight_12_delay_2;
      io_weight_12_delay_4 <= io_weight_12_delay_3;
      io_weight_12_delay_5 <= io_weight_12_delay_4;
      io_weight_12_delay_6 <= io_weight_12_delay_5;
      io_weight_12_delay_7 <= io_weight_12_delay_6;
      io_weight_12_delay_8 <= io_weight_12_delay_7;
      io_weight_12_delay_9 <= io_weight_12_delay_8;
      io_weight_12_delay_10 <= io_weight_12_delay_9;
      io_weight_12_delay_11 <= io_weight_12_delay_10;
      io_weight_12_delay_12 <= io_weight_12_delay_11;
      io_weight_13_delay_1 <= io_weight_13;
      io_weight_13_delay_2 <= io_weight_13_delay_1;
      io_weight_13_delay_3 <= io_weight_13_delay_2;
      io_weight_13_delay_4 <= io_weight_13_delay_3;
      io_weight_13_delay_5 <= io_weight_13_delay_4;
      io_weight_13_delay_6 <= io_weight_13_delay_5;
      io_weight_13_delay_7 <= io_weight_13_delay_6;
      io_weight_13_delay_8 <= io_weight_13_delay_7;
      io_weight_13_delay_9 <= io_weight_13_delay_8;
      io_weight_13_delay_10 <= io_weight_13_delay_9;
      io_weight_13_delay_11 <= io_weight_13_delay_10;
      io_weight_13_delay_12 <= io_weight_13_delay_11;
      io_weight_13_delay_13 <= io_weight_13_delay_12;
      io_weight_14_delay_1 <= io_weight_14;
      io_weight_14_delay_2 <= io_weight_14_delay_1;
      io_weight_14_delay_3 <= io_weight_14_delay_2;
      io_weight_14_delay_4 <= io_weight_14_delay_3;
      io_weight_14_delay_5 <= io_weight_14_delay_4;
      io_weight_14_delay_6 <= io_weight_14_delay_5;
      io_weight_14_delay_7 <= io_weight_14_delay_6;
      io_weight_14_delay_8 <= io_weight_14_delay_7;
      io_weight_14_delay_9 <= io_weight_14_delay_8;
      io_weight_14_delay_10 <= io_weight_14_delay_9;
      io_weight_14_delay_11 <= io_weight_14_delay_10;
      io_weight_14_delay_12 <= io_weight_14_delay_11;
      io_weight_14_delay_13 <= io_weight_14_delay_12;
      io_weight_14_delay_14 <= io_weight_14_delay_13;
      io_weight_15_delay_1 <= io_weight_15;
      io_weight_15_delay_2 <= io_weight_15_delay_1;
      io_weight_15_delay_3 <= io_weight_15_delay_2;
      io_weight_15_delay_4 <= io_weight_15_delay_3;
      io_weight_15_delay_5 <= io_weight_15_delay_4;
      io_weight_15_delay_6 <= io_weight_15_delay_5;
      io_weight_15_delay_7 <= io_weight_15_delay_6;
      io_weight_15_delay_8 <= io_weight_15_delay_7;
      io_weight_15_delay_9 <= io_weight_15_delay_8;
      io_weight_15_delay_10 <= io_weight_15_delay_9;
      io_weight_15_delay_11 <= io_weight_15_delay_10;
      io_weight_15_delay_12 <= io_weight_15_delay_11;
      io_weight_15_delay_13 <= io_weight_15_delay_12;
      io_weight_15_delay_14 <= io_weight_15_delay_13;
      io_weight_15_delay_15 <= io_weight_15_delay_14;
      io_weight_16_delay_1 <= io_weight_16;
      io_weight_16_delay_2 <= io_weight_16_delay_1;
      io_weight_16_delay_3 <= io_weight_16_delay_2;
      io_weight_16_delay_4 <= io_weight_16_delay_3;
      io_weight_16_delay_5 <= io_weight_16_delay_4;
      io_weight_16_delay_6 <= io_weight_16_delay_5;
      io_weight_16_delay_7 <= io_weight_16_delay_6;
      io_weight_16_delay_8 <= io_weight_16_delay_7;
      io_weight_16_delay_9 <= io_weight_16_delay_8;
      io_weight_16_delay_10 <= io_weight_16_delay_9;
      io_weight_16_delay_11 <= io_weight_16_delay_10;
      io_weight_16_delay_12 <= io_weight_16_delay_11;
      io_weight_16_delay_13 <= io_weight_16_delay_12;
      io_weight_16_delay_14 <= io_weight_16_delay_13;
      io_weight_16_delay_15 <= io_weight_16_delay_14;
      io_weight_16_delay_16 <= io_weight_16_delay_15;
      io_weight_17_delay_1 <= io_weight_17;
      io_weight_17_delay_2 <= io_weight_17_delay_1;
      io_weight_17_delay_3 <= io_weight_17_delay_2;
      io_weight_17_delay_4 <= io_weight_17_delay_3;
      io_weight_17_delay_5 <= io_weight_17_delay_4;
      io_weight_17_delay_6 <= io_weight_17_delay_5;
      io_weight_17_delay_7 <= io_weight_17_delay_6;
      io_weight_17_delay_8 <= io_weight_17_delay_7;
      io_weight_17_delay_9 <= io_weight_17_delay_8;
      io_weight_17_delay_10 <= io_weight_17_delay_9;
      io_weight_17_delay_11 <= io_weight_17_delay_10;
      io_weight_17_delay_12 <= io_weight_17_delay_11;
      io_weight_17_delay_13 <= io_weight_17_delay_12;
      io_weight_17_delay_14 <= io_weight_17_delay_13;
      io_weight_17_delay_15 <= io_weight_17_delay_14;
      io_weight_17_delay_16 <= io_weight_17_delay_15;
      io_weight_17_delay_17 <= io_weight_17_delay_16;
      io_weight_18_delay_1 <= io_weight_18;
      io_weight_18_delay_2 <= io_weight_18_delay_1;
      io_weight_18_delay_3 <= io_weight_18_delay_2;
      io_weight_18_delay_4 <= io_weight_18_delay_3;
      io_weight_18_delay_5 <= io_weight_18_delay_4;
      io_weight_18_delay_6 <= io_weight_18_delay_5;
      io_weight_18_delay_7 <= io_weight_18_delay_6;
      io_weight_18_delay_8 <= io_weight_18_delay_7;
      io_weight_18_delay_9 <= io_weight_18_delay_8;
      io_weight_18_delay_10 <= io_weight_18_delay_9;
      io_weight_18_delay_11 <= io_weight_18_delay_10;
      io_weight_18_delay_12 <= io_weight_18_delay_11;
      io_weight_18_delay_13 <= io_weight_18_delay_12;
      io_weight_18_delay_14 <= io_weight_18_delay_13;
      io_weight_18_delay_15 <= io_weight_18_delay_14;
      io_weight_18_delay_16 <= io_weight_18_delay_15;
      io_weight_18_delay_17 <= io_weight_18_delay_16;
      io_weight_18_delay_18 <= io_weight_18_delay_17;
      io_weight_19_delay_1 <= io_weight_19;
      io_weight_19_delay_2 <= io_weight_19_delay_1;
      io_weight_19_delay_3 <= io_weight_19_delay_2;
      io_weight_19_delay_4 <= io_weight_19_delay_3;
      io_weight_19_delay_5 <= io_weight_19_delay_4;
      io_weight_19_delay_6 <= io_weight_19_delay_5;
      io_weight_19_delay_7 <= io_weight_19_delay_6;
      io_weight_19_delay_8 <= io_weight_19_delay_7;
      io_weight_19_delay_9 <= io_weight_19_delay_8;
      io_weight_19_delay_10 <= io_weight_19_delay_9;
      io_weight_19_delay_11 <= io_weight_19_delay_10;
      io_weight_19_delay_12 <= io_weight_19_delay_11;
      io_weight_19_delay_13 <= io_weight_19_delay_12;
      io_weight_19_delay_14 <= io_weight_19_delay_13;
      io_weight_19_delay_15 <= io_weight_19_delay_14;
      io_weight_19_delay_16 <= io_weight_19_delay_15;
      io_weight_19_delay_17 <= io_weight_19_delay_16;
      io_weight_19_delay_18 <= io_weight_19_delay_17;
      io_weight_19_delay_19 <= io_weight_19_delay_18;
      io_weight_20_delay_1 <= io_weight_20;
      io_weight_20_delay_2 <= io_weight_20_delay_1;
      io_weight_20_delay_3 <= io_weight_20_delay_2;
      io_weight_20_delay_4 <= io_weight_20_delay_3;
      io_weight_20_delay_5 <= io_weight_20_delay_4;
      io_weight_20_delay_6 <= io_weight_20_delay_5;
      io_weight_20_delay_7 <= io_weight_20_delay_6;
      io_weight_20_delay_8 <= io_weight_20_delay_7;
      io_weight_20_delay_9 <= io_weight_20_delay_8;
      io_weight_20_delay_10 <= io_weight_20_delay_9;
      io_weight_20_delay_11 <= io_weight_20_delay_10;
      io_weight_20_delay_12 <= io_weight_20_delay_11;
      io_weight_20_delay_13 <= io_weight_20_delay_12;
      io_weight_20_delay_14 <= io_weight_20_delay_13;
      io_weight_20_delay_15 <= io_weight_20_delay_14;
      io_weight_20_delay_16 <= io_weight_20_delay_15;
      io_weight_20_delay_17 <= io_weight_20_delay_16;
      io_weight_20_delay_18 <= io_weight_20_delay_17;
      io_weight_20_delay_19 <= io_weight_20_delay_18;
      io_weight_20_delay_20 <= io_weight_20_delay_19;
      io_weight_21_delay_1 <= io_weight_21;
      io_weight_21_delay_2 <= io_weight_21_delay_1;
      io_weight_21_delay_3 <= io_weight_21_delay_2;
      io_weight_21_delay_4 <= io_weight_21_delay_3;
      io_weight_21_delay_5 <= io_weight_21_delay_4;
      io_weight_21_delay_6 <= io_weight_21_delay_5;
      io_weight_21_delay_7 <= io_weight_21_delay_6;
      io_weight_21_delay_8 <= io_weight_21_delay_7;
      io_weight_21_delay_9 <= io_weight_21_delay_8;
      io_weight_21_delay_10 <= io_weight_21_delay_9;
      io_weight_21_delay_11 <= io_weight_21_delay_10;
      io_weight_21_delay_12 <= io_weight_21_delay_11;
      io_weight_21_delay_13 <= io_weight_21_delay_12;
      io_weight_21_delay_14 <= io_weight_21_delay_13;
      io_weight_21_delay_15 <= io_weight_21_delay_14;
      io_weight_21_delay_16 <= io_weight_21_delay_15;
      io_weight_21_delay_17 <= io_weight_21_delay_16;
      io_weight_21_delay_18 <= io_weight_21_delay_17;
      io_weight_21_delay_19 <= io_weight_21_delay_18;
      io_weight_21_delay_20 <= io_weight_21_delay_19;
      io_weight_21_delay_21 <= io_weight_21_delay_20;
      io_weight_22_delay_1 <= io_weight_22;
      io_weight_22_delay_2 <= io_weight_22_delay_1;
      io_weight_22_delay_3 <= io_weight_22_delay_2;
      io_weight_22_delay_4 <= io_weight_22_delay_3;
      io_weight_22_delay_5 <= io_weight_22_delay_4;
      io_weight_22_delay_6 <= io_weight_22_delay_5;
      io_weight_22_delay_7 <= io_weight_22_delay_6;
      io_weight_22_delay_8 <= io_weight_22_delay_7;
      io_weight_22_delay_9 <= io_weight_22_delay_8;
      io_weight_22_delay_10 <= io_weight_22_delay_9;
      io_weight_22_delay_11 <= io_weight_22_delay_10;
      io_weight_22_delay_12 <= io_weight_22_delay_11;
      io_weight_22_delay_13 <= io_weight_22_delay_12;
      io_weight_22_delay_14 <= io_weight_22_delay_13;
      io_weight_22_delay_15 <= io_weight_22_delay_14;
      io_weight_22_delay_16 <= io_weight_22_delay_15;
      io_weight_22_delay_17 <= io_weight_22_delay_16;
      io_weight_22_delay_18 <= io_weight_22_delay_17;
      io_weight_22_delay_19 <= io_weight_22_delay_18;
      io_weight_22_delay_20 <= io_weight_22_delay_19;
      io_weight_22_delay_21 <= io_weight_22_delay_20;
      io_weight_22_delay_22 <= io_weight_22_delay_21;
      io_weight_23_delay_1 <= io_weight_23;
      io_weight_23_delay_2 <= io_weight_23_delay_1;
      io_weight_23_delay_3 <= io_weight_23_delay_2;
      io_weight_23_delay_4 <= io_weight_23_delay_3;
      io_weight_23_delay_5 <= io_weight_23_delay_4;
      io_weight_23_delay_6 <= io_weight_23_delay_5;
      io_weight_23_delay_7 <= io_weight_23_delay_6;
      io_weight_23_delay_8 <= io_weight_23_delay_7;
      io_weight_23_delay_9 <= io_weight_23_delay_8;
      io_weight_23_delay_10 <= io_weight_23_delay_9;
      io_weight_23_delay_11 <= io_weight_23_delay_10;
      io_weight_23_delay_12 <= io_weight_23_delay_11;
      io_weight_23_delay_13 <= io_weight_23_delay_12;
      io_weight_23_delay_14 <= io_weight_23_delay_13;
      io_weight_23_delay_15 <= io_weight_23_delay_14;
      io_weight_23_delay_16 <= io_weight_23_delay_15;
      io_weight_23_delay_17 <= io_weight_23_delay_16;
      io_weight_23_delay_18 <= io_weight_23_delay_17;
      io_weight_23_delay_19 <= io_weight_23_delay_18;
      io_weight_23_delay_20 <= io_weight_23_delay_19;
      io_weight_23_delay_21 <= io_weight_23_delay_20;
      io_weight_23_delay_22 <= io_weight_23_delay_21;
      io_weight_23_delay_23 <= io_weight_23_delay_22;
      io_weight_24_delay_1 <= io_weight_24;
      io_weight_24_delay_2 <= io_weight_24_delay_1;
      io_weight_24_delay_3 <= io_weight_24_delay_2;
      io_weight_24_delay_4 <= io_weight_24_delay_3;
      io_weight_24_delay_5 <= io_weight_24_delay_4;
      io_weight_24_delay_6 <= io_weight_24_delay_5;
      io_weight_24_delay_7 <= io_weight_24_delay_6;
      io_weight_24_delay_8 <= io_weight_24_delay_7;
      io_weight_24_delay_9 <= io_weight_24_delay_8;
      io_weight_24_delay_10 <= io_weight_24_delay_9;
      io_weight_24_delay_11 <= io_weight_24_delay_10;
      io_weight_24_delay_12 <= io_weight_24_delay_11;
      io_weight_24_delay_13 <= io_weight_24_delay_12;
      io_weight_24_delay_14 <= io_weight_24_delay_13;
      io_weight_24_delay_15 <= io_weight_24_delay_14;
      io_weight_24_delay_16 <= io_weight_24_delay_15;
      io_weight_24_delay_17 <= io_weight_24_delay_16;
      io_weight_24_delay_18 <= io_weight_24_delay_17;
      io_weight_24_delay_19 <= io_weight_24_delay_18;
      io_weight_24_delay_20 <= io_weight_24_delay_19;
      io_weight_24_delay_21 <= io_weight_24_delay_20;
      io_weight_24_delay_22 <= io_weight_24_delay_21;
      io_weight_24_delay_23 <= io_weight_24_delay_22;
      io_weight_24_delay_24 <= io_weight_24_delay_23;
      io_weight_25_delay_1 <= io_weight_25;
      io_weight_25_delay_2 <= io_weight_25_delay_1;
      io_weight_25_delay_3 <= io_weight_25_delay_2;
      io_weight_25_delay_4 <= io_weight_25_delay_3;
      io_weight_25_delay_5 <= io_weight_25_delay_4;
      io_weight_25_delay_6 <= io_weight_25_delay_5;
      io_weight_25_delay_7 <= io_weight_25_delay_6;
      io_weight_25_delay_8 <= io_weight_25_delay_7;
      io_weight_25_delay_9 <= io_weight_25_delay_8;
      io_weight_25_delay_10 <= io_weight_25_delay_9;
      io_weight_25_delay_11 <= io_weight_25_delay_10;
      io_weight_25_delay_12 <= io_weight_25_delay_11;
      io_weight_25_delay_13 <= io_weight_25_delay_12;
      io_weight_25_delay_14 <= io_weight_25_delay_13;
      io_weight_25_delay_15 <= io_weight_25_delay_14;
      io_weight_25_delay_16 <= io_weight_25_delay_15;
      io_weight_25_delay_17 <= io_weight_25_delay_16;
      io_weight_25_delay_18 <= io_weight_25_delay_17;
      io_weight_25_delay_19 <= io_weight_25_delay_18;
      io_weight_25_delay_20 <= io_weight_25_delay_19;
      io_weight_25_delay_21 <= io_weight_25_delay_20;
      io_weight_25_delay_22 <= io_weight_25_delay_21;
      io_weight_25_delay_23 <= io_weight_25_delay_22;
      io_weight_25_delay_24 <= io_weight_25_delay_23;
      io_weight_25_delay_25 <= io_weight_25_delay_24;
      io_weight_26_delay_1 <= io_weight_26;
      io_weight_26_delay_2 <= io_weight_26_delay_1;
      io_weight_26_delay_3 <= io_weight_26_delay_2;
      io_weight_26_delay_4 <= io_weight_26_delay_3;
      io_weight_26_delay_5 <= io_weight_26_delay_4;
      io_weight_26_delay_6 <= io_weight_26_delay_5;
      io_weight_26_delay_7 <= io_weight_26_delay_6;
      io_weight_26_delay_8 <= io_weight_26_delay_7;
      io_weight_26_delay_9 <= io_weight_26_delay_8;
      io_weight_26_delay_10 <= io_weight_26_delay_9;
      io_weight_26_delay_11 <= io_weight_26_delay_10;
      io_weight_26_delay_12 <= io_weight_26_delay_11;
      io_weight_26_delay_13 <= io_weight_26_delay_12;
      io_weight_26_delay_14 <= io_weight_26_delay_13;
      io_weight_26_delay_15 <= io_weight_26_delay_14;
      io_weight_26_delay_16 <= io_weight_26_delay_15;
      io_weight_26_delay_17 <= io_weight_26_delay_16;
      io_weight_26_delay_18 <= io_weight_26_delay_17;
      io_weight_26_delay_19 <= io_weight_26_delay_18;
      io_weight_26_delay_20 <= io_weight_26_delay_19;
      io_weight_26_delay_21 <= io_weight_26_delay_20;
      io_weight_26_delay_22 <= io_weight_26_delay_21;
      io_weight_26_delay_23 <= io_weight_26_delay_22;
      io_weight_26_delay_24 <= io_weight_26_delay_23;
      io_weight_26_delay_25 <= io_weight_26_delay_24;
      io_weight_26_delay_26 <= io_weight_26_delay_25;
      io_weight_27_delay_1 <= io_weight_27;
      io_weight_27_delay_2 <= io_weight_27_delay_1;
      io_weight_27_delay_3 <= io_weight_27_delay_2;
      io_weight_27_delay_4 <= io_weight_27_delay_3;
      io_weight_27_delay_5 <= io_weight_27_delay_4;
      io_weight_27_delay_6 <= io_weight_27_delay_5;
      io_weight_27_delay_7 <= io_weight_27_delay_6;
      io_weight_27_delay_8 <= io_weight_27_delay_7;
      io_weight_27_delay_9 <= io_weight_27_delay_8;
      io_weight_27_delay_10 <= io_weight_27_delay_9;
      io_weight_27_delay_11 <= io_weight_27_delay_10;
      io_weight_27_delay_12 <= io_weight_27_delay_11;
      io_weight_27_delay_13 <= io_weight_27_delay_12;
      io_weight_27_delay_14 <= io_weight_27_delay_13;
      io_weight_27_delay_15 <= io_weight_27_delay_14;
      io_weight_27_delay_16 <= io_weight_27_delay_15;
      io_weight_27_delay_17 <= io_weight_27_delay_16;
      io_weight_27_delay_18 <= io_weight_27_delay_17;
      io_weight_27_delay_19 <= io_weight_27_delay_18;
      io_weight_27_delay_20 <= io_weight_27_delay_19;
      io_weight_27_delay_21 <= io_weight_27_delay_20;
      io_weight_27_delay_22 <= io_weight_27_delay_21;
      io_weight_27_delay_23 <= io_weight_27_delay_22;
      io_weight_27_delay_24 <= io_weight_27_delay_23;
      io_weight_27_delay_25 <= io_weight_27_delay_24;
      io_weight_27_delay_26 <= io_weight_27_delay_25;
      io_weight_27_delay_27 <= io_weight_27_delay_26;
      io_weight_28_delay_1 <= io_weight_28;
      io_weight_28_delay_2 <= io_weight_28_delay_1;
      io_weight_28_delay_3 <= io_weight_28_delay_2;
      io_weight_28_delay_4 <= io_weight_28_delay_3;
      io_weight_28_delay_5 <= io_weight_28_delay_4;
      io_weight_28_delay_6 <= io_weight_28_delay_5;
      io_weight_28_delay_7 <= io_weight_28_delay_6;
      io_weight_28_delay_8 <= io_weight_28_delay_7;
      io_weight_28_delay_9 <= io_weight_28_delay_8;
      io_weight_28_delay_10 <= io_weight_28_delay_9;
      io_weight_28_delay_11 <= io_weight_28_delay_10;
      io_weight_28_delay_12 <= io_weight_28_delay_11;
      io_weight_28_delay_13 <= io_weight_28_delay_12;
      io_weight_28_delay_14 <= io_weight_28_delay_13;
      io_weight_28_delay_15 <= io_weight_28_delay_14;
      io_weight_28_delay_16 <= io_weight_28_delay_15;
      io_weight_28_delay_17 <= io_weight_28_delay_16;
      io_weight_28_delay_18 <= io_weight_28_delay_17;
      io_weight_28_delay_19 <= io_weight_28_delay_18;
      io_weight_28_delay_20 <= io_weight_28_delay_19;
      io_weight_28_delay_21 <= io_weight_28_delay_20;
      io_weight_28_delay_22 <= io_weight_28_delay_21;
      io_weight_28_delay_23 <= io_weight_28_delay_22;
      io_weight_28_delay_24 <= io_weight_28_delay_23;
      io_weight_28_delay_25 <= io_weight_28_delay_24;
      io_weight_28_delay_26 <= io_weight_28_delay_25;
      io_weight_28_delay_27 <= io_weight_28_delay_26;
      io_weight_28_delay_28 <= io_weight_28_delay_27;
      io_weight_29_delay_1 <= io_weight_29;
      io_weight_29_delay_2 <= io_weight_29_delay_1;
      io_weight_29_delay_3 <= io_weight_29_delay_2;
      io_weight_29_delay_4 <= io_weight_29_delay_3;
      io_weight_29_delay_5 <= io_weight_29_delay_4;
      io_weight_29_delay_6 <= io_weight_29_delay_5;
      io_weight_29_delay_7 <= io_weight_29_delay_6;
      io_weight_29_delay_8 <= io_weight_29_delay_7;
      io_weight_29_delay_9 <= io_weight_29_delay_8;
      io_weight_29_delay_10 <= io_weight_29_delay_9;
      io_weight_29_delay_11 <= io_weight_29_delay_10;
      io_weight_29_delay_12 <= io_weight_29_delay_11;
      io_weight_29_delay_13 <= io_weight_29_delay_12;
      io_weight_29_delay_14 <= io_weight_29_delay_13;
      io_weight_29_delay_15 <= io_weight_29_delay_14;
      io_weight_29_delay_16 <= io_weight_29_delay_15;
      io_weight_29_delay_17 <= io_weight_29_delay_16;
      io_weight_29_delay_18 <= io_weight_29_delay_17;
      io_weight_29_delay_19 <= io_weight_29_delay_18;
      io_weight_29_delay_20 <= io_weight_29_delay_19;
      io_weight_29_delay_21 <= io_weight_29_delay_20;
      io_weight_29_delay_22 <= io_weight_29_delay_21;
      io_weight_29_delay_23 <= io_weight_29_delay_22;
      io_weight_29_delay_24 <= io_weight_29_delay_23;
      io_weight_29_delay_25 <= io_weight_29_delay_24;
      io_weight_29_delay_26 <= io_weight_29_delay_25;
      io_weight_29_delay_27 <= io_weight_29_delay_26;
      io_weight_29_delay_28 <= io_weight_29_delay_27;
      io_weight_29_delay_29 <= io_weight_29_delay_28;
      io_weight_30_delay_1 <= io_weight_30;
      io_weight_30_delay_2 <= io_weight_30_delay_1;
      io_weight_30_delay_3 <= io_weight_30_delay_2;
      io_weight_30_delay_4 <= io_weight_30_delay_3;
      io_weight_30_delay_5 <= io_weight_30_delay_4;
      io_weight_30_delay_6 <= io_weight_30_delay_5;
      io_weight_30_delay_7 <= io_weight_30_delay_6;
      io_weight_30_delay_8 <= io_weight_30_delay_7;
      io_weight_30_delay_9 <= io_weight_30_delay_8;
      io_weight_30_delay_10 <= io_weight_30_delay_9;
      io_weight_30_delay_11 <= io_weight_30_delay_10;
      io_weight_30_delay_12 <= io_weight_30_delay_11;
      io_weight_30_delay_13 <= io_weight_30_delay_12;
      io_weight_30_delay_14 <= io_weight_30_delay_13;
      io_weight_30_delay_15 <= io_weight_30_delay_14;
      io_weight_30_delay_16 <= io_weight_30_delay_15;
      io_weight_30_delay_17 <= io_weight_30_delay_16;
      io_weight_30_delay_18 <= io_weight_30_delay_17;
      io_weight_30_delay_19 <= io_weight_30_delay_18;
      io_weight_30_delay_20 <= io_weight_30_delay_19;
      io_weight_30_delay_21 <= io_weight_30_delay_20;
      io_weight_30_delay_22 <= io_weight_30_delay_21;
      io_weight_30_delay_23 <= io_weight_30_delay_22;
      io_weight_30_delay_24 <= io_weight_30_delay_23;
      io_weight_30_delay_25 <= io_weight_30_delay_24;
      io_weight_30_delay_26 <= io_weight_30_delay_25;
      io_weight_30_delay_27 <= io_weight_30_delay_26;
      io_weight_30_delay_28 <= io_weight_30_delay_27;
      io_weight_30_delay_29 <= io_weight_30_delay_28;
      io_weight_30_delay_30 <= io_weight_30_delay_29;
      io_weight_31_delay_1 <= io_weight_31;
      io_weight_31_delay_2 <= io_weight_31_delay_1;
      io_weight_31_delay_3 <= io_weight_31_delay_2;
      io_weight_31_delay_4 <= io_weight_31_delay_3;
      io_weight_31_delay_5 <= io_weight_31_delay_4;
      io_weight_31_delay_6 <= io_weight_31_delay_5;
      io_weight_31_delay_7 <= io_weight_31_delay_6;
      io_weight_31_delay_8 <= io_weight_31_delay_7;
      io_weight_31_delay_9 <= io_weight_31_delay_8;
      io_weight_31_delay_10 <= io_weight_31_delay_9;
      io_weight_31_delay_11 <= io_weight_31_delay_10;
      io_weight_31_delay_12 <= io_weight_31_delay_11;
      io_weight_31_delay_13 <= io_weight_31_delay_12;
      io_weight_31_delay_14 <= io_weight_31_delay_13;
      io_weight_31_delay_15 <= io_weight_31_delay_14;
      io_weight_31_delay_16 <= io_weight_31_delay_15;
      io_weight_31_delay_17 <= io_weight_31_delay_16;
      io_weight_31_delay_18 <= io_weight_31_delay_17;
      io_weight_31_delay_19 <= io_weight_31_delay_18;
      io_weight_31_delay_20 <= io_weight_31_delay_19;
      io_weight_31_delay_21 <= io_weight_31_delay_20;
      io_weight_31_delay_22 <= io_weight_31_delay_21;
      io_weight_31_delay_23 <= io_weight_31_delay_22;
      io_weight_31_delay_24 <= io_weight_31_delay_23;
      io_weight_31_delay_25 <= io_weight_31_delay_24;
      io_weight_31_delay_26 <= io_weight_31_delay_25;
      io_weight_31_delay_27 <= io_weight_31_delay_26;
      io_weight_31_delay_28 <= io_weight_31_delay_27;
      io_weight_31_delay_29 <= io_weight_31_delay_28;
      io_weight_31_delay_30 <= io_weight_31_delay_29;
      io_weight_31_delay_31 <= io_weight_31_delay_30;
      toplevel_mac_0_31_io_macOut_delay_1 <= mac_0_31_io_macOut;
      toplevel_mac_0_31_io_macOut_delay_2 <= toplevel_mac_0_31_io_macOut_delay_1;
      toplevel_mac_0_31_io_macOut_delay_3 <= toplevel_mac_0_31_io_macOut_delay_2;
      toplevel_mac_0_31_io_macOut_delay_4 <= toplevel_mac_0_31_io_macOut_delay_3;
      toplevel_mac_0_31_io_macOut_delay_5 <= toplevel_mac_0_31_io_macOut_delay_4;
      toplevel_mac_0_31_io_macOut_delay_6 <= toplevel_mac_0_31_io_macOut_delay_5;
      toplevel_mac_0_31_io_macOut_delay_7 <= toplevel_mac_0_31_io_macOut_delay_6;
      toplevel_mac_0_31_io_macOut_delay_8 <= toplevel_mac_0_31_io_macOut_delay_7;
      toplevel_mac_0_31_io_macOut_delay_9 <= toplevel_mac_0_31_io_macOut_delay_8;
      toplevel_mac_0_31_io_macOut_delay_10 <= toplevel_mac_0_31_io_macOut_delay_9;
      toplevel_mac_0_31_io_macOut_delay_11 <= toplevel_mac_0_31_io_macOut_delay_10;
      toplevel_mac_0_31_io_macOut_delay_12 <= toplevel_mac_0_31_io_macOut_delay_11;
      toplevel_mac_0_31_io_macOut_delay_13 <= toplevel_mac_0_31_io_macOut_delay_12;
      toplevel_mac_0_31_io_macOut_delay_14 <= toplevel_mac_0_31_io_macOut_delay_13;
      toplevel_mac_0_31_io_macOut_delay_15 <= toplevel_mac_0_31_io_macOut_delay_14;
      toplevel_mac_0_31_io_macOut_delay_16 <= toplevel_mac_0_31_io_macOut_delay_15;
      toplevel_mac_0_31_io_macOut_delay_17 <= toplevel_mac_0_31_io_macOut_delay_16;
      toplevel_mac_0_31_io_macOut_delay_18 <= toplevel_mac_0_31_io_macOut_delay_17;
      toplevel_mac_0_31_io_macOut_delay_19 <= toplevel_mac_0_31_io_macOut_delay_18;
      toplevel_mac_0_31_io_macOut_delay_20 <= toplevel_mac_0_31_io_macOut_delay_19;
      toplevel_mac_0_31_io_macOut_delay_21 <= toplevel_mac_0_31_io_macOut_delay_20;
      toplevel_mac_0_31_io_macOut_delay_22 <= toplevel_mac_0_31_io_macOut_delay_21;
      toplevel_mac_0_31_io_macOut_delay_23 <= toplevel_mac_0_31_io_macOut_delay_22;
      toplevel_mac_0_31_io_macOut_delay_24 <= toplevel_mac_0_31_io_macOut_delay_23;
      toplevel_mac_0_31_io_macOut_delay_25 <= toplevel_mac_0_31_io_macOut_delay_24;
      toplevel_mac_0_31_io_macOut_delay_26 <= toplevel_mac_0_31_io_macOut_delay_25;
      toplevel_mac_0_31_io_macOut_delay_27 <= toplevel_mac_0_31_io_macOut_delay_26;
      toplevel_mac_0_31_io_macOut_delay_28 <= toplevel_mac_0_31_io_macOut_delay_27;
      toplevel_mac_0_31_io_macOut_delay_29 <= toplevel_mac_0_31_io_macOut_delay_28;
      toplevel_mac_0_31_io_macOut_delay_30 <= toplevel_mac_0_31_io_macOut_delay_29;
      toplevel_mac_0_31_io_macOut_delay_31 <= toplevel_mac_0_31_io_macOut_delay_30;
      toplevel_mac_1_31_io_macOut_delay_1 <= mac_1_31_io_macOut;
      toplevel_mac_1_31_io_macOut_delay_2 <= toplevel_mac_1_31_io_macOut_delay_1;
      toplevel_mac_1_31_io_macOut_delay_3 <= toplevel_mac_1_31_io_macOut_delay_2;
      toplevel_mac_1_31_io_macOut_delay_4 <= toplevel_mac_1_31_io_macOut_delay_3;
      toplevel_mac_1_31_io_macOut_delay_5 <= toplevel_mac_1_31_io_macOut_delay_4;
      toplevel_mac_1_31_io_macOut_delay_6 <= toplevel_mac_1_31_io_macOut_delay_5;
      toplevel_mac_1_31_io_macOut_delay_7 <= toplevel_mac_1_31_io_macOut_delay_6;
      toplevel_mac_1_31_io_macOut_delay_8 <= toplevel_mac_1_31_io_macOut_delay_7;
      toplevel_mac_1_31_io_macOut_delay_9 <= toplevel_mac_1_31_io_macOut_delay_8;
      toplevel_mac_1_31_io_macOut_delay_10 <= toplevel_mac_1_31_io_macOut_delay_9;
      toplevel_mac_1_31_io_macOut_delay_11 <= toplevel_mac_1_31_io_macOut_delay_10;
      toplevel_mac_1_31_io_macOut_delay_12 <= toplevel_mac_1_31_io_macOut_delay_11;
      toplevel_mac_1_31_io_macOut_delay_13 <= toplevel_mac_1_31_io_macOut_delay_12;
      toplevel_mac_1_31_io_macOut_delay_14 <= toplevel_mac_1_31_io_macOut_delay_13;
      toplevel_mac_1_31_io_macOut_delay_15 <= toplevel_mac_1_31_io_macOut_delay_14;
      toplevel_mac_1_31_io_macOut_delay_16 <= toplevel_mac_1_31_io_macOut_delay_15;
      toplevel_mac_1_31_io_macOut_delay_17 <= toplevel_mac_1_31_io_macOut_delay_16;
      toplevel_mac_1_31_io_macOut_delay_18 <= toplevel_mac_1_31_io_macOut_delay_17;
      toplevel_mac_1_31_io_macOut_delay_19 <= toplevel_mac_1_31_io_macOut_delay_18;
      toplevel_mac_1_31_io_macOut_delay_20 <= toplevel_mac_1_31_io_macOut_delay_19;
      toplevel_mac_1_31_io_macOut_delay_21 <= toplevel_mac_1_31_io_macOut_delay_20;
      toplevel_mac_1_31_io_macOut_delay_22 <= toplevel_mac_1_31_io_macOut_delay_21;
      toplevel_mac_1_31_io_macOut_delay_23 <= toplevel_mac_1_31_io_macOut_delay_22;
      toplevel_mac_1_31_io_macOut_delay_24 <= toplevel_mac_1_31_io_macOut_delay_23;
      toplevel_mac_1_31_io_macOut_delay_25 <= toplevel_mac_1_31_io_macOut_delay_24;
      toplevel_mac_1_31_io_macOut_delay_26 <= toplevel_mac_1_31_io_macOut_delay_25;
      toplevel_mac_1_31_io_macOut_delay_27 <= toplevel_mac_1_31_io_macOut_delay_26;
      toplevel_mac_1_31_io_macOut_delay_28 <= toplevel_mac_1_31_io_macOut_delay_27;
      toplevel_mac_1_31_io_macOut_delay_29 <= toplevel_mac_1_31_io_macOut_delay_28;
      toplevel_mac_1_31_io_macOut_delay_30 <= toplevel_mac_1_31_io_macOut_delay_29;
      toplevel_mac_2_31_io_macOut_delay_1 <= mac_2_31_io_macOut;
      toplevel_mac_2_31_io_macOut_delay_2 <= toplevel_mac_2_31_io_macOut_delay_1;
      toplevel_mac_2_31_io_macOut_delay_3 <= toplevel_mac_2_31_io_macOut_delay_2;
      toplevel_mac_2_31_io_macOut_delay_4 <= toplevel_mac_2_31_io_macOut_delay_3;
      toplevel_mac_2_31_io_macOut_delay_5 <= toplevel_mac_2_31_io_macOut_delay_4;
      toplevel_mac_2_31_io_macOut_delay_6 <= toplevel_mac_2_31_io_macOut_delay_5;
      toplevel_mac_2_31_io_macOut_delay_7 <= toplevel_mac_2_31_io_macOut_delay_6;
      toplevel_mac_2_31_io_macOut_delay_8 <= toplevel_mac_2_31_io_macOut_delay_7;
      toplevel_mac_2_31_io_macOut_delay_9 <= toplevel_mac_2_31_io_macOut_delay_8;
      toplevel_mac_2_31_io_macOut_delay_10 <= toplevel_mac_2_31_io_macOut_delay_9;
      toplevel_mac_2_31_io_macOut_delay_11 <= toplevel_mac_2_31_io_macOut_delay_10;
      toplevel_mac_2_31_io_macOut_delay_12 <= toplevel_mac_2_31_io_macOut_delay_11;
      toplevel_mac_2_31_io_macOut_delay_13 <= toplevel_mac_2_31_io_macOut_delay_12;
      toplevel_mac_2_31_io_macOut_delay_14 <= toplevel_mac_2_31_io_macOut_delay_13;
      toplevel_mac_2_31_io_macOut_delay_15 <= toplevel_mac_2_31_io_macOut_delay_14;
      toplevel_mac_2_31_io_macOut_delay_16 <= toplevel_mac_2_31_io_macOut_delay_15;
      toplevel_mac_2_31_io_macOut_delay_17 <= toplevel_mac_2_31_io_macOut_delay_16;
      toplevel_mac_2_31_io_macOut_delay_18 <= toplevel_mac_2_31_io_macOut_delay_17;
      toplevel_mac_2_31_io_macOut_delay_19 <= toplevel_mac_2_31_io_macOut_delay_18;
      toplevel_mac_2_31_io_macOut_delay_20 <= toplevel_mac_2_31_io_macOut_delay_19;
      toplevel_mac_2_31_io_macOut_delay_21 <= toplevel_mac_2_31_io_macOut_delay_20;
      toplevel_mac_2_31_io_macOut_delay_22 <= toplevel_mac_2_31_io_macOut_delay_21;
      toplevel_mac_2_31_io_macOut_delay_23 <= toplevel_mac_2_31_io_macOut_delay_22;
      toplevel_mac_2_31_io_macOut_delay_24 <= toplevel_mac_2_31_io_macOut_delay_23;
      toplevel_mac_2_31_io_macOut_delay_25 <= toplevel_mac_2_31_io_macOut_delay_24;
      toplevel_mac_2_31_io_macOut_delay_26 <= toplevel_mac_2_31_io_macOut_delay_25;
      toplevel_mac_2_31_io_macOut_delay_27 <= toplevel_mac_2_31_io_macOut_delay_26;
      toplevel_mac_2_31_io_macOut_delay_28 <= toplevel_mac_2_31_io_macOut_delay_27;
      toplevel_mac_2_31_io_macOut_delay_29 <= toplevel_mac_2_31_io_macOut_delay_28;
      toplevel_mac_3_31_io_macOut_delay_1 <= mac_3_31_io_macOut;
      toplevel_mac_3_31_io_macOut_delay_2 <= toplevel_mac_3_31_io_macOut_delay_1;
      toplevel_mac_3_31_io_macOut_delay_3 <= toplevel_mac_3_31_io_macOut_delay_2;
      toplevel_mac_3_31_io_macOut_delay_4 <= toplevel_mac_3_31_io_macOut_delay_3;
      toplevel_mac_3_31_io_macOut_delay_5 <= toplevel_mac_3_31_io_macOut_delay_4;
      toplevel_mac_3_31_io_macOut_delay_6 <= toplevel_mac_3_31_io_macOut_delay_5;
      toplevel_mac_3_31_io_macOut_delay_7 <= toplevel_mac_3_31_io_macOut_delay_6;
      toplevel_mac_3_31_io_macOut_delay_8 <= toplevel_mac_3_31_io_macOut_delay_7;
      toplevel_mac_3_31_io_macOut_delay_9 <= toplevel_mac_3_31_io_macOut_delay_8;
      toplevel_mac_3_31_io_macOut_delay_10 <= toplevel_mac_3_31_io_macOut_delay_9;
      toplevel_mac_3_31_io_macOut_delay_11 <= toplevel_mac_3_31_io_macOut_delay_10;
      toplevel_mac_3_31_io_macOut_delay_12 <= toplevel_mac_3_31_io_macOut_delay_11;
      toplevel_mac_3_31_io_macOut_delay_13 <= toplevel_mac_3_31_io_macOut_delay_12;
      toplevel_mac_3_31_io_macOut_delay_14 <= toplevel_mac_3_31_io_macOut_delay_13;
      toplevel_mac_3_31_io_macOut_delay_15 <= toplevel_mac_3_31_io_macOut_delay_14;
      toplevel_mac_3_31_io_macOut_delay_16 <= toplevel_mac_3_31_io_macOut_delay_15;
      toplevel_mac_3_31_io_macOut_delay_17 <= toplevel_mac_3_31_io_macOut_delay_16;
      toplevel_mac_3_31_io_macOut_delay_18 <= toplevel_mac_3_31_io_macOut_delay_17;
      toplevel_mac_3_31_io_macOut_delay_19 <= toplevel_mac_3_31_io_macOut_delay_18;
      toplevel_mac_3_31_io_macOut_delay_20 <= toplevel_mac_3_31_io_macOut_delay_19;
      toplevel_mac_3_31_io_macOut_delay_21 <= toplevel_mac_3_31_io_macOut_delay_20;
      toplevel_mac_3_31_io_macOut_delay_22 <= toplevel_mac_3_31_io_macOut_delay_21;
      toplevel_mac_3_31_io_macOut_delay_23 <= toplevel_mac_3_31_io_macOut_delay_22;
      toplevel_mac_3_31_io_macOut_delay_24 <= toplevel_mac_3_31_io_macOut_delay_23;
      toplevel_mac_3_31_io_macOut_delay_25 <= toplevel_mac_3_31_io_macOut_delay_24;
      toplevel_mac_3_31_io_macOut_delay_26 <= toplevel_mac_3_31_io_macOut_delay_25;
      toplevel_mac_3_31_io_macOut_delay_27 <= toplevel_mac_3_31_io_macOut_delay_26;
      toplevel_mac_3_31_io_macOut_delay_28 <= toplevel_mac_3_31_io_macOut_delay_27;
      toplevel_mac_4_31_io_macOut_delay_1 <= mac_4_31_io_macOut;
      toplevel_mac_4_31_io_macOut_delay_2 <= toplevel_mac_4_31_io_macOut_delay_1;
      toplevel_mac_4_31_io_macOut_delay_3 <= toplevel_mac_4_31_io_macOut_delay_2;
      toplevel_mac_4_31_io_macOut_delay_4 <= toplevel_mac_4_31_io_macOut_delay_3;
      toplevel_mac_4_31_io_macOut_delay_5 <= toplevel_mac_4_31_io_macOut_delay_4;
      toplevel_mac_4_31_io_macOut_delay_6 <= toplevel_mac_4_31_io_macOut_delay_5;
      toplevel_mac_4_31_io_macOut_delay_7 <= toplevel_mac_4_31_io_macOut_delay_6;
      toplevel_mac_4_31_io_macOut_delay_8 <= toplevel_mac_4_31_io_macOut_delay_7;
      toplevel_mac_4_31_io_macOut_delay_9 <= toplevel_mac_4_31_io_macOut_delay_8;
      toplevel_mac_4_31_io_macOut_delay_10 <= toplevel_mac_4_31_io_macOut_delay_9;
      toplevel_mac_4_31_io_macOut_delay_11 <= toplevel_mac_4_31_io_macOut_delay_10;
      toplevel_mac_4_31_io_macOut_delay_12 <= toplevel_mac_4_31_io_macOut_delay_11;
      toplevel_mac_4_31_io_macOut_delay_13 <= toplevel_mac_4_31_io_macOut_delay_12;
      toplevel_mac_4_31_io_macOut_delay_14 <= toplevel_mac_4_31_io_macOut_delay_13;
      toplevel_mac_4_31_io_macOut_delay_15 <= toplevel_mac_4_31_io_macOut_delay_14;
      toplevel_mac_4_31_io_macOut_delay_16 <= toplevel_mac_4_31_io_macOut_delay_15;
      toplevel_mac_4_31_io_macOut_delay_17 <= toplevel_mac_4_31_io_macOut_delay_16;
      toplevel_mac_4_31_io_macOut_delay_18 <= toplevel_mac_4_31_io_macOut_delay_17;
      toplevel_mac_4_31_io_macOut_delay_19 <= toplevel_mac_4_31_io_macOut_delay_18;
      toplevel_mac_4_31_io_macOut_delay_20 <= toplevel_mac_4_31_io_macOut_delay_19;
      toplevel_mac_4_31_io_macOut_delay_21 <= toplevel_mac_4_31_io_macOut_delay_20;
      toplevel_mac_4_31_io_macOut_delay_22 <= toplevel_mac_4_31_io_macOut_delay_21;
      toplevel_mac_4_31_io_macOut_delay_23 <= toplevel_mac_4_31_io_macOut_delay_22;
      toplevel_mac_4_31_io_macOut_delay_24 <= toplevel_mac_4_31_io_macOut_delay_23;
      toplevel_mac_4_31_io_macOut_delay_25 <= toplevel_mac_4_31_io_macOut_delay_24;
      toplevel_mac_4_31_io_macOut_delay_26 <= toplevel_mac_4_31_io_macOut_delay_25;
      toplevel_mac_4_31_io_macOut_delay_27 <= toplevel_mac_4_31_io_macOut_delay_26;
      toplevel_mac_5_31_io_macOut_delay_1 <= mac_5_31_io_macOut;
      toplevel_mac_5_31_io_macOut_delay_2 <= toplevel_mac_5_31_io_macOut_delay_1;
      toplevel_mac_5_31_io_macOut_delay_3 <= toplevel_mac_5_31_io_macOut_delay_2;
      toplevel_mac_5_31_io_macOut_delay_4 <= toplevel_mac_5_31_io_macOut_delay_3;
      toplevel_mac_5_31_io_macOut_delay_5 <= toplevel_mac_5_31_io_macOut_delay_4;
      toplevel_mac_5_31_io_macOut_delay_6 <= toplevel_mac_5_31_io_macOut_delay_5;
      toplevel_mac_5_31_io_macOut_delay_7 <= toplevel_mac_5_31_io_macOut_delay_6;
      toplevel_mac_5_31_io_macOut_delay_8 <= toplevel_mac_5_31_io_macOut_delay_7;
      toplevel_mac_5_31_io_macOut_delay_9 <= toplevel_mac_5_31_io_macOut_delay_8;
      toplevel_mac_5_31_io_macOut_delay_10 <= toplevel_mac_5_31_io_macOut_delay_9;
      toplevel_mac_5_31_io_macOut_delay_11 <= toplevel_mac_5_31_io_macOut_delay_10;
      toplevel_mac_5_31_io_macOut_delay_12 <= toplevel_mac_5_31_io_macOut_delay_11;
      toplevel_mac_5_31_io_macOut_delay_13 <= toplevel_mac_5_31_io_macOut_delay_12;
      toplevel_mac_5_31_io_macOut_delay_14 <= toplevel_mac_5_31_io_macOut_delay_13;
      toplevel_mac_5_31_io_macOut_delay_15 <= toplevel_mac_5_31_io_macOut_delay_14;
      toplevel_mac_5_31_io_macOut_delay_16 <= toplevel_mac_5_31_io_macOut_delay_15;
      toplevel_mac_5_31_io_macOut_delay_17 <= toplevel_mac_5_31_io_macOut_delay_16;
      toplevel_mac_5_31_io_macOut_delay_18 <= toplevel_mac_5_31_io_macOut_delay_17;
      toplevel_mac_5_31_io_macOut_delay_19 <= toplevel_mac_5_31_io_macOut_delay_18;
      toplevel_mac_5_31_io_macOut_delay_20 <= toplevel_mac_5_31_io_macOut_delay_19;
      toplevel_mac_5_31_io_macOut_delay_21 <= toplevel_mac_5_31_io_macOut_delay_20;
      toplevel_mac_5_31_io_macOut_delay_22 <= toplevel_mac_5_31_io_macOut_delay_21;
      toplevel_mac_5_31_io_macOut_delay_23 <= toplevel_mac_5_31_io_macOut_delay_22;
      toplevel_mac_5_31_io_macOut_delay_24 <= toplevel_mac_5_31_io_macOut_delay_23;
      toplevel_mac_5_31_io_macOut_delay_25 <= toplevel_mac_5_31_io_macOut_delay_24;
      toplevel_mac_5_31_io_macOut_delay_26 <= toplevel_mac_5_31_io_macOut_delay_25;
      toplevel_mac_6_31_io_macOut_delay_1 <= mac_6_31_io_macOut;
      toplevel_mac_6_31_io_macOut_delay_2 <= toplevel_mac_6_31_io_macOut_delay_1;
      toplevel_mac_6_31_io_macOut_delay_3 <= toplevel_mac_6_31_io_macOut_delay_2;
      toplevel_mac_6_31_io_macOut_delay_4 <= toplevel_mac_6_31_io_macOut_delay_3;
      toplevel_mac_6_31_io_macOut_delay_5 <= toplevel_mac_6_31_io_macOut_delay_4;
      toplevel_mac_6_31_io_macOut_delay_6 <= toplevel_mac_6_31_io_macOut_delay_5;
      toplevel_mac_6_31_io_macOut_delay_7 <= toplevel_mac_6_31_io_macOut_delay_6;
      toplevel_mac_6_31_io_macOut_delay_8 <= toplevel_mac_6_31_io_macOut_delay_7;
      toplevel_mac_6_31_io_macOut_delay_9 <= toplevel_mac_6_31_io_macOut_delay_8;
      toplevel_mac_6_31_io_macOut_delay_10 <= toplevel_mac_6_31_io_macOut_delay_9;
      toplevel_mac_6_31_io_macOut_delay_11 <= toplevel_mac_6_31_io_macOut_delay_10;
      toplevel_mac_6_31_io_macOut_delay_12 <= toplevel_mac_6_31_io_macOut_delay_11;
      toplevel_mac_6_31_io_macOut_delay_13 <= toplevel_mac_6_31_io_macOut_delay_12;
      toplevel_mac_6_31_io_macOut_delay_14 <= toplevel_mac_6_31_io_macOut_delay_13;
      toplevel_mac_6_31_io_macOut_delay_15 <= toplevel_mac_6_31_io_macOut_delay_14;
      toplevel_mac_6_31_io_macOut_delay_16 <= toplevel_mac_6_31_io_macOut_delay_15;
      toplevel_mac_6_31_io_macOut_delay_17 <= toplevel_mac_6_31_io_macOut_delay_16;
      toplevel_mac_6_31_io_macOut_delay_18 <= toplevel_mac_6_31_io_macOut_delay_17;
      toplevel_mac_6_31_io_macOut_delay_19 <= toplevel_mac_6_31_io_macOut_delay_18;
      toplevel_mac_6_31_io_macOut_delay_20 <= toplevel_mac_6_31_io_macOut_delay_19;
      toplevel_mac_6_31_io_macOut_delay_21 <= toplevel_mac_6_31_io_macOut_delay_20;
      toplevel_mac_6_31_io_macOut_delay_22 <= toplevel_mac_6_31_io_macOut_delay_21;
      toplevel_mac_6_31_io_macOut_delay_23 <= toplevel_mac_6_31_io_macOut_delay_22;
      toplevel_mac_6_31_io_macOut_delay_24 <= toplevel_mac_6_31_io_macOut_delay_23;
      toplevel_mac_6_31_io_macOut_delay_25 <= toplevel_mac_6_31_io_macOut_delay_24;
      toplevel_mac_7_31_io_macOut_delay_1 <= mac_7_31_io_macOut;
      toplevel_mac_7_31_io_macOut_delay_2 <= toplevel_mac_7_31_io_macOut_delay_1;
      toplevel_mac_7_31_io_macOut_delay_3 <= toplevel_mac_7_31_io_macOut_delay_2;
      toplevel_mac_7_31_io_macOut_delay_4 <= toplevel_mac_7_31_io_macOut_delay_3;
      toplevel_mac_7_31_io_macOut_delay_5 <= toplevel_mac_7_31_io_macOut_delay_4;
      toplevel_mac_7_31_io_macOut_delay_6 <= toplevel_mac_7_31_io_macOut_delay_5;
      toplevel_mac_7_31_io_macOut_delay_7 <= toplevel_mac_7_31_io_macOut_delay_6;
      toplevel_mac_7_31_io_macOut_delay_8 <= toplevel_mac_7_31_io_macOut_delay_7;
      toplevel_mac_7_31_io_macOut_delay_9 <= toplevel_mac_7_31_io_macOut_delay_8;
      toplevel_mac_7_31_io_macOut_delay_10 <= toplevel_mac_7_31_io_macOut_delay_9;
      toplevel_mac_7_31_io_macOut_delay_11 <= toplevel_mac_7_31_io_macOut_delay_10;
      toplevel_mac_7_31_io_macOut_delay_12 <= toplevel_mac_7_31_io_macOut_delay_11;
      toplevel_mac_7_31_io_macOut_delay_13 <= toplevel_mac_7_31_io_macOut_delay_12;
      toplevel_mac_7_31_io_macOut_delay_14 <= toplevel_mac_7_31_io_macOut_delay_13;
      toplevel_mac_7_31_io_macOut_delay_15 <= toplevel_mac_7_31_io_macOut_delay_14;
      toplevel_mac_7_31_io_macOut_delay_16 <= toplevel_mac_7_31_io_macOut_delay_15;
      toplevel_mac_7_31_io_macOut_delay_17 <= toplevel_mac_7_31_io_macOut_delay_16;
      toplevel_mac_7_31_io_macOut_delay_18 <= toplevel_mac_7_31_io_macOut_delay_17;
      toplevel_mac_7_31_io_macOut_delay_19 <= toplevel_mac_7_31_io_macOut_delay_18;
      toplevel_mac_7_31_io_macOut_delay_20 <= toplevel_mac_7_31_io_macOut_delay_19;
      toplevel_mac_7_31_io_macOut_delay_21 <= toplevel_mac_7_31_io_macOut_delay_20;
      toplevel_mac_7_31_io_macOut_delay_22 <= toplevel_mac_7_31_io_macOut_delay_21;
      toplevel_mac_7_31_io_macOut_delay_23 <= toplevel_mac_7_31_io_macOut_delay_22;
      toplevel_mac_7_31_io_macOut_delay_24 <= toplevel_mac_7_31_io_macOut_delay_23;
      toplevel_mac_8_31_io_macOut_delay_1 <= mac_8_31_io_macOut;
      toplevel_mac_8_31_io_macOut_delay_2 <= toplevel_mac_8_31_io_macOut_delay_1;
      toplevel_mac_8_31_io_macOut_delay_3 <= toplevel_mac_8_31_io_macOut_delay_2;
      toplevel_mac_8_31_io_macOut_delay_4 <= toplevel_mac_8_31_io_macOut_delay_3;
      toplevel_mac_8_31_io_macOut_delay_5 <= toplevel_mac_8_31_io_macOut_delay_4;
      toplevel_mac_8_31_io_macOut_delay_6 <= toplevel_mac_8_31_io_macOut_delay_5;
      toplevel_mac_8_31_io_macOut_delay_7 <= toplevel_mac_8_31_io_macOut_delay_6;
      toplevel_mac_8_31_io_macOut_delay_8 <= toplevel_mac_8_31_io_macOut_delay_7;
      toplevel_mac_8_31_io_macOut_delay_9 <= toplevel_mac_8_31_io_macOut_delay_8;
      toplevel_mac_8_31_io_macOut_delay_10 <= toplevel_mac_8_31_io_macOut_delay_9;
      toplevel_mac_8_31_io_macOut_delay_11 <= toplevel_mac_8_31_io_macOut_delay_10;
      toplevel_mac_8_31_io_macOut_delay_12 <= toplevel_mac_8_31_io_macOut_delay_11;
      toplevel_mac_8_31_io_macOut_delay_13 <= toplevel_mac_8_31_io_macOut_delay_12;
      toplevel_mac_8_31_io_macOut_delay_14 <= toplevel_mac_8_31_io_macOut_delay_13;
      toplevel_mac_8_31_io_macOut_delay_15 <= toplevel_mac_8_31_io_macOut_delay_14;
      toplevel_mac_8_31_io_macOut_delay_16 <= toplevel_mac_8_31_io_macOut_delay_15;
      toplevel_mac_8_31_io_macOut_delay_17 <= toplevel_mac_8_31_io_macOut_delay_16;
      toplevel_mac_8_31_io_macOut_delay_18 <= toplevel_mac_8_31_io_macOut_delay_17;
      toplevel_mac_8_31_io_macOut_delay_19 <= toplevel_mac_8_31_io_macOut_delay_18;
      toplevel_mac_8_31_io_macOut_delay_20 <= toplevel_mac_8_31_io_macOut_delay_19;
      toplevel_mac_8_31_io_macOut_delay_21 <= toplevel_mac_8_31_io_macOut_delay_20;
      toplevel_mac_8_31_io_macOut_delay_22 <= toplevel_mac_8_31_io_macOut_delay_21;
      toplevel_mac_8_31_io_macOut_delay_23 <= toplevel_mac_8_31_io_macOut_delay_22;
      toplevel_mac_9_31_io_macOut_delay_1 <= mac_9_31_io_macOut;
      toplevel_mac_9_31_io_macOut_delay_2 <= toplevel_mac_9_31_io_macOut_delay_1;
      toplevel_mac_9_31_io_macOut_delay_3 <= toplevel_mac_9_31_io_macOut_delay_2;
      toplevel_mac_9_31_io_macOut_delay_4 <= toplevel_mac_9_31_io_macOut_delay_3;
      toplevel_mac_9_31_io_macOut_delay_5 <= toplevel_mac_9_31_io_macOut_delay_4;
      toplevel_mac_9_31_io_macOut_delay_6 <= toplevel_mac_9_31_io_macOut_delay_5;
      toplevel_mac_9_31_io_macOut_delay_7 <= toplevel_mac_9_31_io_macOut_delay_6;
      toplevel_mac_9_31_io_macOut_delay_8 <= toplevel_mac_9_31_io_macOut_delay_7;
      toplevel_mac_9_31_io_macOut_delay_9 <= toplevel_mac_9_31_io_macOut_delay_8;
      toplevel_mac_9_31_io_macOut_delay_10 <= toplevel_mac_9_31_io_macOut_delay_9;
      toplevel_mac_9_31_io_macOut_delay_11 <= toplevel_mac_9_31_io_macOut_delay_10;
      toplevel_mac_9_31_io_macOut_delay_12 <= toplevel_mac_9_31_io_macOut_delay_11;
      toplevel_mac_9_31_io_macOut_delay_13 <= toplevel_mac_9_31_io_macOut_delay_12;
      toplevel_mac_9_31_io_macOut_delay_14 <= toplevel_mac_9_31_io_macOut_delay_13;
      toplevel_mac_9_31_io_macOut_delay_15 <= toplevel_mac_9_31_io_macOut_delay_14;
      toplevel_mac_9_31_io_macOut_delay_16 <= toplevel_mac_9_31_io_macOut_delay_15;
      toplevel_mac_9_31_io_macOut_delay_17 <= toplevel_mac_9_31_io_macOut_delay_16;
      toplevel_mac_9_31_io_macOut_delay_18 <= toplevel_mac_9_31_io_macOut_delay_17;
      toplevel_mac_9_31_io_macOut_delay_19 <= toplevel_mac_9_31_io_macOut_delay_18;
      toplevel_mac_9_31_io_macOut_delay_20 <= toplevel_mac_9_31_io_macOut_delay_19;
      toplevel_mac_9_31_io_macOut_delay_21 <= toplevel_mac_9_31_io_macOut_delay_20;
      toplevel_mac_9_31_io_macOut_delay_22 <= toplevel_mac_9_31_io_macOut_delay_21;
      toplevel_mac_10_31_io_macOut_delay_1 <= mac_10_31_io_macOut;
      toplevel_mac_10_31_io_macOut_delay_2 <= toplevel_mac_10_31_io_macOut_delay_1;
      toplevel_mac_10_31_io_macOut_delay_3 <= toplevel_mac_10_31_io_macOut_delay_2;
      toplevel_mac_10_31_io_macOut_delay_4 <= toplevel_mac_10_31_io_macOut_delay_3;
      toplevel_mac_10_31_io_macOut_delay_5 <= toplevel_mac_10_31_io_macOut_delay_4;
      toplevel_mac_10_31_io_macOut_delay_6 <= toplevel_mac_10_31_io_macOut_delay_5;
      toplevel_mac_10_31_io_macOut_delay_7 <= toplevel_mac_10_31_io_macOut_delay_6;
      toplevel_mac_10_31_io_macOut_delay_8 <= toplevel_mac_10_31_io_macOut_delay_7;
      toplevel_mac_10_31_io_macOut_delay_9 <= toplevel_mac_10_31_io_macOut_delay_8;
      toplevel_mac_10_31_io_macOut_delay_10 <= toplevel_mac_10_31_io_macOut_delay_9;
      toplevel_mac_10_31_io_macOut_delay_11 <= toplevel_mac_10_31_io_macOut_delay_10;
      toplevel_mac_10_31_io_macOut_delay_12 <= toplevel_mac_10_31_io_macOut_delay_11;
      toplevel_mac_10_31_io_macOut_delay_13 <= toplevel_mac_10_31_io_macOut_delay_12;
      toplevel_mac_10_31_io_macOut_delay_14 <= toplevel_mac_10_31_io_macOut_delay_13;
      toplevel_mac_10_31_io_macOut_delay_15 <= toplevel_mac_10_31_io_macOut_delay_14;
      toplevel_mac_10_31_io_macOut_delay_16 <= toplevel_mac_10_31_io_macOut_delay_15;
      toplevel_mac_10_31_io_macOut_delay_17 <= toplevel_mac_10_31_io_macOut_delay_16;
      toplevel_mac_10_31_io_macOut_delay_18 <= toplevel_mac_10_31_io_macOut_delay_17;
      toplevel_mac_10_31_io_macOut_delay_19 <= toplevel_mac_10_31_io_macOut_delay_18;
      toplevel_mac_10_31_io_macOut_delay_20 <= toplevel_mac_10_31_io_macOut_delay_19;
      toplevel_mac_10_31_io_macOut_delay_21 <= toplevel_mac_10_31_io_macOut_delay_20;
      toplevel_mac_11_31_io_macOut_delay_1 <= mac_11_31_io_macOut;
      toplevel_mac_11_31_io_macOut_delay_2 <= toplevel_mac_11_31_io_macOut_delay_1;
      toplevel_mac_11_31_io_macOut_delay_3 <= toplevel_mac_11_31_io_macOut_delay_2;
      toplevel_mac_11_31_io_macOut_delay_4 <= toplevel_mac_11_31_io_macOut_delay_3;
      toplevel_mac_11_31_io_macOut_delay_5 <= toplevel_mac_11_31_io_macOut_delay_4;
      toplevel_mac_11_31_io_macOut_delay_6 <= toplevel_mac_11_31_io_macOut_delay_5;
      toplevel_mac_11_31_io_macOut_delay_7 <= toplevel_mac_11_31_io_macOut_delay_6;
      toplevel_mac_11_31_io_macOut_delay_8 <= toplevel_mac_11_31_io_macOut_delay_7;
      toplevel_mac_11_31_io_macOut_delay_9 <= toplevel_mac_11_31_io_macOut_delay_8;
      toplevel_mac_11_31_io_macOut_delay_10 <= toplevel_mac_11_31_io_macOut_delay_9;
      toplevel_mac_11_31_io_macOut_delay_11 <= toplevel_mac_11_31_io_macOut_delay_10;
      toplevel_mac_11_31_io_macOut_delay_12 <= toplevel_mac_11_31_io_macOut_delay_11;
      toplevel_mac_11_31_io_macOut_delay_13 <= toplevel_mac_11_31_io_macOut_delay_12;
      toplevel_mac_11_31_io_macOut_delay_14 <= toplevel_mac_11_31_io_macOut_delay_13;
      toplevel_mac_11_31_io_macOut_delay_15 <= toplevel_mac_11_31_io_macOut_delay_14;
      toplevel_mac_11_31_io_macOut_delay_16 <= toplevel_mac_11_31_io_macOut_delay_15;
      toplevel_mac_11_31_io_macOut_delay_17 <= toplevel_mac_11_31_io_macOut_delay_16;
      toplevel_mac_11_31_io_macOut_delay_18 <= toplevel_mac_11_31_io_macOut_delay_17;
      toplevel_mac_11_31_io_macOut_delay_19 <= toplevel_mac_11_31_io_macOut_delay_18;
      toplevel_mac_11_31_io_macOut_delay_20 <= toplevel_mac_11_31_io_macOut_delay_19;
      toplevel_mac_12_31_io_macOut_delay_1 <= mac_12_31_io_macOut;
      toplevel_mac_12_31_io_macOut_delay_2 <= toplevel_mac_12_31_io_macOut_delay_1;
      toplevel_mac_12_31_io_macOut_delay_3 <= toplevel_mac_12_31_io_macOut_delay_2;
      toplevel_mac_12_31_io_macOut_delay_4 <= toplevel_mac_12_31_io_macOut_delay_3;
      toplevel_mac_12_31_io_macOut_delay_5 <= toplevel_mac_12_31_io_macOut_delay_4;
      toplevel_mac_12_31_io_macOut_delay_6 <= toplevel_mac_12_31_io_macOut_delay_5;
      toplevel_mac_12_31_io_macOut_delay_7 <= toplevel_mac_12_31_io_macOut_delay_6;
      toplevel_mac_12_31_io_macOut_delay_8 <= toplevel_mac_12_31_io_macOut_delay_7;
      toplevel_mac_12_31_io_macOut_delay_9 <= toplevel_mac_12_31_io_macOut_delay_8;
      toplevel_mac_12_31_io_macOut_delay_10 <= toplevel_mac_12_31_io_macOut_delay_9;
      toplevel_mac_12_31_io_macOut_delay_11 <= toplevel_mac_12_31_io_macOut_delay_10;
      toplevel_mac_12_31_io_macOut_delay_12 <= toplevel_mac_12_31_io_macOut_delay_11;
      toplevel_mac_12_31_io_macOut_delay_13 <= toplevel_mac_12_31_io_macOut_delay_12;
      toplevel_mac_12_31_io_macOut_delay_14 <= toplevel_mac_12_31_io_macOut_delay_13;
      toplevel_mac_12_31_io_macOut_delay_15 <= toplevel_mac_12_31_io_macOut_delay_14;
      toplevel_mac_12_31_io_macOut_delay_16 <= toplevel_mac_12_31_io_macOut_delay_15;
      toplevel_mac_12_31_io_macOut_delay_17 <= toplevel_mac_12_31_io_macOut_delay_16;
      toplevel_mac_12_31_io_macOut_delay_18 <= toplevel_mac_12_31_io_macOut_delay_17;
      toplevel_mac_12_31_io_macOut_delay_19 <= toplevel_mac_12_31_io_macOut_delay_18;
      toplevel_mac_13_31_io_macOut_delay_1 <= mac_13_31_io_macOut;
      toplevel_mac_13_31_io_macOut_delay_2 <= toplevel_mac_13_31_io_macOut_delay_1;
      toplevel_mac_13_31_io_macOut_delay_3 <= toplevel_mac_13_31_io_macOut_delay_2;
      toplevel_mac_13_31_io_macOut_delay_4 <= toplevel_mac_13_31_io_macOut_delay_3;
      toplevel_mac_13_31_io_macOut_delay_5 <= toplevel_mac_13_31_io_macOut_delay_4;
      toplevel_mac_13_31_io_macOut_delay_6 <= toplevel_mac_13_31_io_macOut_delay_5;
      toplevel_mac_13_31_io_macOut_delay_7 <= toplevel_mac_13_31_io_macOut_delay_6;
      toplevel_mac_13_31_io_macOut_delay_8 <= toplevel_mac_13_31_io_macOut_delay_7;
      toplevel_mac_13_31_io_macOut_delay_9 <= toplevel_mac_13_31_io_macOut_delay_8;
      toplevel_mac_13_31_io_macOut_delay_10 <= toplevel_mac_13_31_io_macOut_delay_9;
      toplevel_mac_13_31_io_macOut_delay_11 <= toplevel_mac_13_31_io_macOut_delay_10;
      toplevel_mac_13_31_io_macOut_delay_12 <= toplevel_mac_13_31_io_macOut_delay_11;
      toplevel_mac_13_31_io_macOut_delay_13 <= toplevel_mac_13_31_io_macOut_delay_12;
      toplevel_mac_13_31_io_macOut_delay_14 <= toplevel_mac_13_31_io_macOut_delay_13;
      toplevel_mac_13_31_io_macOut_delay_15 <= toplevel_mac_13_31_io_macOut_delay_14;
      toplevel_mac_13_31_io_macOut_delay_16 <= toplevel_mac_13_31_io_macOut_delay_15;
      toplevel_mac_13_31_io_macOut_delay_17 <= toplevel_mac_13_31_io_macOut_delay_16;
      toplevel_mac_13_31_io_macOut_delay_18 <= toplevel_mac_13_31_io_macOut_delay_17;
      toplevel_mac_14_31_io_macOut_delay_1 <= mac_14_31_io_macOut;
      toplevel_mac_14_31_io_macOut_delay_2 <= toplevel_mac_14_31_io_macOut_delay_1;
      toplevel_mac_14_31_io_macOut_delay_3 <= toplevel_mac_14_31_io_macOut_delay_2;
      toplevel_mac_14_31_io_macOut_delay_4 <= toplevel_mac_14_31_io_macOut_delay_3;
      toplevel_mac_14_31_io_macOut_delay_5 <= toplevel_mac_14_31_io_macOut_delay_4;
      toplevel_mac_14_31_io_macOut_delay_6 <= toplevel_mac_14_31_io_macOut_delay_5;
      toplevel_mac_14_31_io_macOut_delay_7 <= toplevel_mac_14_31_io_macOut_delay_6;
      toplevel_mac_14_31_io_macOut_delay_8 <= toplevel_mac_14_31_io_macOut_delay_7;
      toplevel_mac_14_31_io_macOut_delay_9 <= toplevel_mac_14_31_io_macOut_delay_8;
      toplevel_mac_14_31_io_macOut_delay_10 <= toplevel_mac_14_31_io_macOut_delay_9;
      toplevel_mac_14_31_io_macOut_delay_11 <= toplevel_mac_14_31_io_macOut_delay_10;
      toplevel_mac_14_31_io_macOut_delay_12 <= toplevel_mac_14_31_io_macOut_delay_11;
      toplevel_mac_14_31_io_macOut_delay_13 <= toplevel_mac_14_31_io_macOut_delay_12;
      toplevel_mac_14_31_io_macOut_delay_14 <= toplevel_mac_14_31_io_macOut_delay_13;
      toplevel_mac_14_31_io_macOut_delay_15 <= toplevel_mac_14_31_io_macOut_delay_14;
      toplevel_mac_14_31_io_macOut_delay_16 <= toplevel_mac_14_31_io_macOut_delay_15;
      toplevel_mac_14_31_io_macOut_delay_17 <= toplevel_mac_14_31_io_macOut_delay_16;
      toplevel_mac_15_31_io_macOut_delay_1 <= mac_15_31_io_macOut;
      toplevel_mac_15_31_io_macOut_delay_2 <= toplevel_mac_15_31_io_macOut_delay_1;
      toplevel_mac_15_31_io_macOut_delay_3 <= toplevel_mac_15_31_io_macOut_delay_2;
      toplevel_mac_15_31_io_macOut_delay_4 <= toplevel_mac_15_31_io_macOut_delay_3;
      toplevel_mac_15_31_io_macOut_delay_5 <= toplevel_mac_15_31_io_macOut_delay_4;
      toplevel_mac_15_31_io_macOut_delay_6 <= toplevel_mac_15_31_io_macOut_delay_5;
      toplevel_mac_15_31_io_macOut_delay_7 <= toplevel_mac_15_31_io_macOut_delay_6;
      toplevel_mac_15_31_io_macOut_delay_8 <= toplevel_mac_15_31_io_macOut_delay_7;
      toplevel_mac_15_31_io_macOut_delay_9 <= toplevel_mac_15_31_io_macOut_delay_8;
      toplevel_mac_15_31_io_macOut_delay_10 <= toplevel_mac_15_31_io_macOut_delay_9;
      toplevel_mac_15_31_io_macOut_delay_11 <= toplevel_mac_15_31_io_macOut_delay_10;
      toplevel_mac_15_31_io_macOut_delay_12 <= toplevel_mac_15_31_io_macOut_delay_11;
      toplevel_mac_15_31_io_macOut_delay_13 <= toplevel_mac_15_31_io_macOut_delay_12;
      toplevel_mac_15_31_io_macOut_delay_14 <= toplevel_mac_15_31_io_macOut_delay_13;
      toplevel_mac_15_31_io_macOut_delay_15 <= toplevel_mac_15_31_io_macOut_delay_14;
      toplevel_mac_15_31_io_macOut_delay_16 <= toplevel_mac_15_31_io_macOut_delay_15;
      toplevel_mac_16_31_io_macOut_delay_1 <= mac_16_31_io_macOut;
      toplevel_mac_16_31_io_macOut_delay_2 <= toplevel_mac_16_31_io_macOut_delay_1;
      toplevel_mac_16_31_io_macOut_delay_3 <= toplevel_mac_16_31_io_macOut_delay_2;
      toplevel_mac_16_31_io_macOut_delay_4 <= toplevel_mac_16_31_io_macOut_delay_3;
      toplevel_mac_16_31_io_macOut_delay_5 <= toplevel_mac_16_31_io_macOut_delay_4;
      toplevel_mac_16_31_io_macOut_delay_6 <= toplevel_mac_16_31_io_macOut_delay_5;
      toplevel_mac_16_31_io_macOut_delay_7 <= toplevel_mac_16_31_io_macOut_delay_6;
      toplevel_mac_16_31_io_macOut_delay_8 <= toplevel_mac_16_31_io_macOut_delay_7;
      toplevel_mac_16_31_io_macOut_delay_9 <= toplevel_mac_16_31_io_macOut_delay_8;
      toplevel_mac_16_31_io_macOut_delay_10 <= toplevel_mac_16_31_io_macOut_delay_9;
      toplevel_mac_16_31_io_macOut_delay_11 <= toplevel_mac_16_31_io_macOut_delay_10;
      toplevel_mac_16_31_io_macOut_delay_12 <= toplevel_mac_16_31_io_macOut_delay_11;
      toplevel_mac_16_31_io_macOut_delay_13 <= toplevel_mac_16_31_io_macOut_delay_12;
      toplevel_mac_16_31_io_macOut_delay_14 <= toplevel_mac_16_31_io_macOut_delay_13;
      toplevel_mac_16_31_io_macOut_delay_15 <= toplevel_mac_16_31_io_macOut_delay_14;
      toplevel_mac_17_31_io_macOut_delay_1 <= mac_17_31_io_macOut;
      toplevel_mac_17_31_io_macOut_delay_2 <= toplevel_mac_17_31_io_macOut_delay_1;
      toplevel_mac_17_31_io_macOut_delay_3 <= toplevel_mac_17_31_io_macOut_delay_2;
      toplevel_mac_17_31_io_macOut_delay_4 <= toplevel_mac_17_31_io_macOut_delay_3;
      toplevel_mac_17_31_io_macOut_delay_5 <= toplevel_mac_17_31_io_macOut_delay_4;
      toplevel_mac_17_31_io_macOut_delay_6 <= toplevel_mac_17_31_io_macOut_delay_5;
      toplevel_mac_17_31_io_macOut_delay_7 <= toplevel_mac_17_31_io_macOut_delay_6;
      toplevel_mac_17_31_io_macOut_delay_8 <= toplevel_mac_17_31_io_macOut_delay_7;
      toplevel_mac_17_31_io_macOut_delay_9 <= toplevel_mac_17_31_io_macOut_delay_8;
      toplevel_mac_17_31_io_macOut_delay_10 <= toplevel_mac_17_31_io_macOut_delay_9;
      toplevel_mac_17_31_io_macOut_delay_11 <= toplevel_mac_17_31_io_macOut_delay_10;
      toplevel_mac_17_31_io_macOut_delay_12 <= toplevel_mac_17_31_io_macOut_delay_11;
      toplevel_mac_17_31_io_macOut_delay_13 <= toplevel_mac_17_31_io_macOut_delay_12;
      toplevel_mac_17_31_io_macOut_delay_14 <= toplevel_mac_17_31_io_macOut_delay_13;
      toplevel_mac_18_31_io_macOut_delay_1 <= mac_18_31_io_macOut;
      toplevel_mac_18_31_io_macOut_delay_2 <= toplevel_mac_18_31_io_macOut_delay_1;
      toplevel_mac_18_31_io_macOut_delay_3 <= toplevel_mac_18_31_io_macOut_delay_2;
      toplevel_mac_18_31_io_macOut_delay_4 <= toplevel_mac_18_31_io_macOut_delay_3;
      toplevel_mac_18_31_io_macOut_delay_5 <= toplevel_mac_18_31_io_macOut_delay_4;
      toplevel_mac_18_31_io_macOut_delay_6 <= toplevel_mac_18_31_io_macOut_delay_5;
      toplevel_mac_18_31_io_macOut_delay_7 <= toplevel_mac_18_31_io_macOut_delay_6;
      toplevel_mac_18_31_io_macOut_delay_8 <= toplevel_mac_18_31_io_macOut_delay_7;
      toplevel_mac_18_31_io_macOut_delay_9 <= toplevel_mac_18_31_io_macOut_delay_8;
      toplevel_mac_18_31_io_macOut_delay_10 <= toplevel_mac_18_31_io_macOut_delay_9;
      toplevel_mac_18_31_io_macOut_delay_11 <= toplevel_mac_18_31_io_macOut_delay_10;
      toplevel_mac_18_31_io_macOut_delay_12 <= toplevel_mac_18_31_io_macOut_delay_11;
      toplevel_mac_18_31_io_macOut_delay_13 <= toplevel_mac_18_31_io_macOut_delay_12;
      toplevel_mac_19_31_io_macOut_delay_1 <= mac_19_31_io_macOut;
      toplevel_mac_19_31_io_macOut_delay_2 <= toplevel_mac_19_31_io_macOut_delay_1;
      toplevel_mac_19_31_io_macOut_delay_3 <= toplevel_mac_19_31_io_macOut_delay_2;
      toplevel_mac_19_31_io_macOut_delay_4 <= toplevel_mac_19_31_io_macOut_delay_3;
      toplevel_mac_19_31_io_macOut_delay_5 <= toplevel_mac_19_31_io_macOut_delay_4;
      toplevel_mac_19_31_io_macOut_delay_6 <= toplevel_mac_19_31_io_macOut_delay_5;
      toplevel_mac_19_31_io_macOut_delay_7 <= toplevel_mac_19_31_io_macOut_delay_6;
      toplevel_mac_19_31_io_macOut_delay_8 <= toplevel_mac_19_31_io_macOut_delay_7;
      toplevel_mac_19_31_io_macOut_delay_9 <= toplevel_mac_19_31_io_macOut_delay_8;
      toplevel_mac_19_31_io_macOut_delay_10 <= toplevel_mac_19_31_io_macOut_delay_9;
      toplevel_mac_19_31_io_macOut_delay_11 <= toplevel_mac_19_31_io_macOut_delay_10;
      toplevel_mac_19_31_io_macOut_delay_12 <= toplevel_mac_19_31_io_macOut_delay_11;
      toplevel_mac_20_31_io_macOut_delay_1 <= mac_20_31_io_macOut;
      toplevel_mac_20_31_io_macOut_delay_2 <= toplevel_mac_20_31_io_macOut_delay_1;
      toplevel_mac_20_31_io_macOut_delay_3 <= toplevel_mac_20_31_io_macOut_delay_2;
      toplevel_mac_20_31_io_macOut_delay_4 <= toplevel_mac_20_31_io_macOut_delay_3;
      toplevel_mac_20_31_io_macOut_delay_5 <= toplevel_mac_20_31_io_macOut_delay_4;
      toplevel_mac_20_31_io_macOut_delay_6 <= toplevel_mac_20_31_io_macOut_delay_5;
      toplevel_mac_20_31_io_macOut_delay_7 <= toplevel_mac_20_31_io_macOut_delay_6;
      toplevel_mac_20_31_io_macOut_delay_8 <= toplevel_mac_20_31_io_macOut_delay_7;
      toplevel_mac_20_31_io_macOut_delay_9 <= toplevel_mac_20_31_io_macOut_delay_8;
      toplevel_mac_20_31_io_macOut_delay_10 <= toplevel_mac_20_31_io_macOut_delay_9;
      toplevel_mac_20_31_io_macOut_delay_11 <= toplevel_mac_20_31_io_macOut_delay_10;
      toplevel_mac_21_31_io_macOut_delay_1 <= mac_21_31_io_macOut;
      toplevel_mac_21_31_io_macOut_delay_2 <= toplevel_mac_21_31_io_macOut_delay_1;
      toplevel_mac_21_31_io_macOut_delay_3 <= toplevel_mac_21_31_io_macOut_delay_2;
      toplevel_mac_21_31_io_macOut_delay_4 <= toplevel_mac_21_31_io_macOut_delay_3;
      toplevel_mac_21_31_io_macOut_delay_5 <= toplevel_mac_21_31_io_macOut_delay_4;
      toplevel_mac_21_31_io_macOut_delay_6 <= toplevel_mac_21_31_io_macOut_delay_5;
      toplevel_mac_21_31_io_macOut_delay_7 <= toplevel_mac_21_31_io_macOut_delay_6;
      toplevel_mac_21_31_io_macOut_delay_8 <= toplevel_mac_21_31_io_macOut_delay_7;
      toplevel_mac_21_31_io_macOut_delay_9 <= toplevel_mac_21_31_io_macOut_delay_8;
      toplevel_mac_21_31_io_macOut_delay_10 <= toplevel_mac_21_31_io_macOut_delay_9;
      toplevel_mac_22_31_io_macOut_delay_1 <= mac_22_31_io_macOut;
      toplevel_mac_22_31_io_macOut_delay_2 <= toplevel_mac_22_31_io_macOut_delay_1;
      toplevel_mac_22_31_io_macOut_delay_3 <= toplevel_mac_22_31_io_macOut_delay_2;
      toplevel_mac_22_31_io_macOut_delay_4 <= toplevel_mac_22_31_io_macOut_delay_3;
      toplevel_mac_22_31_io_macOut_delay_5 <= toplevel_mac_22_31_io_macOut_delay_4;
      toplevel_mac_22_31_io_macOut_delay_6 <= toplevel_mac_22_31_io_macOut_delay_5;
      toplevel_mac_22_31_io_macOut_delay_7 <= toplevel_mac_22_31_io_macOut_delay_6;
      toplevel_mac_22_31_io_macOut_delay_8 <= toplevel_mac_22_31_io_macOut_delay_7;
      toplevel_mac_22_31_io_macOut_delay_9 <= toplevel_mac_22_31_io_macOut_delay_8;
      toplevel_mac_23_31_io_macOut_delay_1 <= mac_23_31_io_macOut;
      toplevel_mac_23_31_io_macOut_delay_2 <= toplevel_mac_23_31_io_macOut_delay_1;
      toplevel_mac_23_31_io_macOut_delay_3 <= toplevel_mac_23_31_io_macOut_delay_2;
      toplevel_mac_23_31_io_macOut_delay_4 <= toplevel_mac_23_31_io_macOut_delay_3;
      toplevel_mac_23_31_io_macOut_delay_5 <= toplevel_mac_23_31_io_macOut_delay_4;
      toplevel_mac_23_31_io_macOut_delay_6 <= toplevel_mac_23_31_io_macOut_delay_5;
      toplevel_mac_23_31_io_macOut_delay_7 <= toplevel_mac_23_31_io_macOut_delay_6;
      toplevel_mac_23_31_io_macOut_delay_8 <= toplevel_mac_23_31_io_macOut_delay_7;
      toplevel_mac_24_31_io_macOut_delay_1 <= mac_24_31_io_macOut;
      toplevel_mac_24_31_io_macOut_delay_2 <= toplevel_mac_24_31_io_macOut_delay_1;
      toplevel_mac_24_31_io_macOut_delay_3 <= toplevel_mac_24_31_io_macOut_delay_2;
      toplevel_mac_24_31_io_macOut_delay_4 <= toplevel_mac_24_31_io_macOut_delay_3;
      toplevel_mac_24_31_io_macOut_delay_5 <= toplevel_mac_24_31_io_macOut_delay_4;
      toplevel_mac_24_31_io_macOut_delay_6 <= toplevel_mac_24_31_io_macOut_delay_5;
      toplevel_mac_24_31_io_macOut_delay_7 <= toplevel_mac_24_31_io_macOut_delay_6;
      toplevel_mac_25_31_io_macOut_delay_1 <= mac_25_31_io_macOut;
      toplevel_mac_25_31_io_macOut_delay_2 <= toplevel_mac_25_31_io_macOut_delay_1;
      toplevel_mac_25_31_io_macOut_delay_3 <= toplevel_mac_25_31_io_macOut_delay_2;
      toplevel_mac_25_31_io_macOut_delay_4 <= toplevel_mac_25_31_io_macOut_delay_3;
      toplevel_mac_25_31_io_macOut_delay_5 <= toplevel_mac_25_31_io_macOut_delay_4;
      toplevel_mac_25_31_io_macOut_delay_6 <= toplevel_mac_25_31_io_macOut_delay_5;
      toplevel_mac_26_31_io_macOut_delay_1 <= mac_26_31_io_macOut;
      toplevel_mac_26_31_io_macOut_delay_2 <= toplevel_mac_26_31_io_macOut_delay_1;
      toplevel_mac_26_31_io_macOut_delay_3 <= toplevel_mac_26_31_io_macOut_delay_2;
      toplevel_mac_26_31_io_macOut_delay_4 <= toplevel_mac_26_31_io_macOut_delay_3;
      toplevel_mac_26_31_io_macOut_delay_5 <= toplevel_mac_26_31_io_macOut_delay_4;
      toplevel_mac_27_31_io_macOut_delay_1 <= mac_27_31_io_macOut;
      toplevel_mac_27_31_io_macOut_delay_2 <= toplevel_mac_27_31_io_macOut_delay_1;
      toplevel_mac_27_31_io_macOut_delay_3 <= toplevel_mac_27_31_io_macOut_delay_2;
      toplevel_mac_27_31_io_macOut_delay_4 <= toplevel_mac_27_31_io_macOut_delay_3;
      toplevel_mac_28_31_io_macOut_delay_1 <= mac_28_31_io_macOut;
      toplevel_mac_28_31_io_macOut_delay_2 <= toplevel_mac_28_31_io_macOut_delay_1;
      toplevel_mac_28_31_io_macOut_delay_3 <= toplevel_mac_28_31_io_macOut_delay_2;
      toplevel_mac_29_31_io_macOut_delay_1 <= mac_29_31_io_macOut;
      toplevel_mac_29_31_io_macOut_delay_2 <= toplevel_mac_29_31_io_macOut_delay_1;
      toplevel_mac_30_31_io_macOut_delay_1 <= mac_30_31_io_macOut;
    end
  end


endmodule

module MAC_1023 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_31_inner_macOut;
  wire       [15:0]   _zz__zz__31_31_inner_macOut_1;
  wire       [15:0]   _zz__31_31_inner_macOut_1;
  wire       [15:0]   _zz__31_31_inner_macOut_2;
  reg        [7:0]    _31_31_inner_activation;
  reg        [7:0]    _31_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_31_inner_macOut;

  assign _zz__zz__31_31_inner_macOut = ($signed(io_mulInput) * $signed(_31_31_inner_activation));
  assign _zz__zz__31_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_31_inner_macOut)) ? 16'h007f : _zz__31_31_inner_macOut_2);
  assign _zz__31_31_inner_macOut_2 = (($signed(_zz__31_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_31_inner_activation;
    end else begin
      io_macOut = _31_31_inner_macOut;
    end
  end

  assign _zz__31_31_inner_macOut = ($signed(_zz__zz__31_31_inner_macOut) + $signed(_zz__zz__31_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_31_inner_activation <= 8'h00;
      _31_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_31_inner_activation <= io_addInput;
      end else begin
        _31_31_inner_macOut <= _zz__31_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1022 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_30_inner_macOut;
  wire       [15:0]   _zz__zz__31_30_inner_macOut_1;
  wire       [15:0]   _zz__31_30_inner_macOut_1;
  wire       [15:0]   _zz__31_30_inner_macOut_2;
  reg        [7:0]    _31_30_inner_activation;
  reg        [7:0]    _31_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_30_inner_macOut;

  assign _zz__zz__31_30_inner_macOut = ($signed(io_mulInput) * $signed(_31_30_inner_activation));
  assign _zz__zz__31_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_30_inner_macOut)) ? 16'h007f : _zz__31_30_inner_macOut_2);
  assign _zz__31_30_inner_macOut_2 = (($signed(_zz__31_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_30_inner_activation;
    end else begin
      io_macOut = _31_30_inner_macOut;
    end
  end

  assign _zz__31_30_inner_macOut = ($signed(_zz__zz__31_30_inner_macOut) + $signed(_zz__zz__31_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_30_inner_activation <= 8'h00;
      _31_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_30_inner_activation <= io_addInput;
      end else begin
        _31_30_inner_macOut <= _zz__31_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1021 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_29_inner_macOut;
  wire       [15:0]   _zz__zz__31_29_inner_macOut_1;
  wire       [15:0]   _zz__31_29_inner_macOut_1;
  wire       [15:0]   _zz__31_29_inner_macOut_2;
  reg        [7:0]    _31_29_inner_activation;
  reg        [7:0]    _31_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_29_inner_macOut;

  assign _zz__zz__31_29_inner_macOut = ($signed(io_mulInput) * $signed(_31_29_inner_activation));
  assign _zz__zz__31_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_29_inner_macOut)) ? 16'h007f : _zz__31_29_inner_macOut_2);
  assign _zz__31_29_inner_macOut_2 = (($signed(_zz__31_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_29_inner_activation;
    end else begin
      io_macOut = _31_29_inner_macOut;
    end
  end

  assign _zz__31_29_inner_macOut = ($signed(_zz__zz__31_29_inner_macOut) + $signed(_zz__zz__31_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_29_inner_activation <= 8'h00;
      _31_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_29_inner_activation <= io_addInput;
      end else begin
        _31_29_inner_macOut <= _zz__31_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1020 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_28_inner_macOut;
  wire       [15:0]   _zz__zz__31_28_inner_macOut_1;
  wire       [15:0]   _zz__31_28_inner_macOut_1;
  wire       [15:0]   _zz__31_28_inner_macOut_2;
  reg        [7:0]    _31_28_inner_activation;
  reg        [7:0]    _31_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_28_inner_macOut;

  assign _zz__zz__31_28_inner_macOut = ($signed(io_mulInput) * $signed(_31_28_inner_activation));
  assign _zz__zz__31_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_28_inner_macOut)) ? 16'h007f : _zz__31_28_inner_macOut_2);
  assign _zz__31_28_inner_macOut_2 = (($signed(_zz__31_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_28_inner_activation;
    end else begin
      io_macOut = _31_28_inner_macOut;
    end
  end

  assign _zz__31_28_inner_macOut = ($signed(_zz__zz__31_28_inner_macOut) + $signed(_zz__zz__31_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_28_inner_activation <= 8'h00;
      _31_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_28_inner_activation <= io_addInput;
      end else begin
        _31_28_inner_macOut <= _zz__31_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1019 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_27_inner_macOut;
  wire       [15:0]   _zz__zz__31_27_inner_macOut_1;
  wire       [15:0]   _zz__31_27_inner_macOut_1;
  wire       [15:0]   _zz__31_27_inner_macOut_2;
  reg        [7:0]    _31_27_inner_activation;
  reg        [7:0]    _31_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_27_inner_macOut;

  assign _zz__zz__31_27_inner_macOut = ($signed(io_mulInput) * $signed(_31_27_inner_activation));
  assign _zz__zz__31_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_27_inner_macOut)) ? 16'h007f : _zz__31_27_inner_macOut_2);
  assign _zz__31_27_inner_macOut_2 = (($signed(_zz__31_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_27_inner_activation;
    end else begin
      io_macOut = _31_27_inner_macOut;
    end
  end

  assign _zz__31_27_inner_macOut = ($signed(_zz__zz__31_27_inner_macOut) + $signed(_zz__zz__31_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_27_inner_activation <= 8'h00;
      _31_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_27_inner_activation <= io_addInput;
      end else begin
        _31_27_inner_macOut <= _zz__31_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1018 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_26_inner_macOut;
  wire       [15:0]   _zz__zz__31_26_inner_macOut_1;
  wire       [15:0]   _zz__31_26_inner_macOut_1;
  wire       [15:0]   _zz__31_26_inner_macOut_2;
  reg        [7:0]    _31_26_inner_activation;
  reg        [7:0]    _31_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_26_inner_macOut;

  assign _zz__zz__31_26_inner_macOut = ($signed(io_mulInput) * $signed(_31_26_inner_activation));
  assign _zz__zz__31_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_26_inner_macOut)) ? 16'h007f : _zz__31_26_inner_macOut_2);
  assign _zz__31_26_inner_macOut_2 = (($signed(_zz__31_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_26_inner_activation;
    end else begin
      io_macOut = _31_26_inner_macOut;
    end
  end

  assign _zz__31_26_inner_macOut = ($signed(_zz__zz__31_26_inner_macOut) + $signed(_zz__zz__31_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_26_inner_activation <= 8'h00;
      _31_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_26_inner_activation <= io_addInput;
      end else begin
        _31_26_inner_macOut <= _zz__31_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1017 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_25_inner_macOut;
  wire       [15:0]   _zz__zz__31_25_inner_macOut_1;
  wire       [15:0]   _zz__31_25_inner_macOut_1;
  wire       [15:0]   _zz__31_25_inner_macOut_2;
  reg        [7:0]    _31_25_inner_activation;
  reg        [7:0]    _31_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_25_inner_macOut;

  assign _zz__zz__31_25_inner_macOut = ($signed(io_mulInput) * $signed(_31_25_inner_activation));
  assign _zz__zz__31_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_25_inner_macOut)) ? 16'h007f : _zz__31_25_inner_macOut_2);
  assign _zz__31_25_inner_macOut_2 = (($signed(_zz__31_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_25_inner_activation;
    end else begin
      io_macOut = _31_25_inner_macOut;
    end
  end

  assign _zz__31_25_inner_macOut = ($signed(_zz__zz__31_25_inner_macOut) + $signed(_zz__zz__31_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_25_inner_activation <= 8'h00;
      _31_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_25_inner_activation <= io_addInput;
      end else begin
        _31_25_inner_macOut <= _zz__31_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1016 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_24_inner_macOut;
  wire       [15:0]   _zz__zz__31_24_inner_macOut_1;
  wire       [15:0]   _zz__31_24_inner_macOut_1;
  wire       [15:0]   _zz__31_24_inner_macOut_2;
  reg        [7:0]    _31_24_inner_activation;
  reg        [7:0]    _31_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_24_inner_macOut;

  assign _zz__zz__31_24_inner_macOut = ($signed(io_mulInput) * $signed(_31_24_inner_activation));
  assign _zz__zz__31_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_24_inner_macOut)) ? 16'h007f : _zz__31_24_inner_macOut_2);
  assign _zz__31_24_inner_macOut_2 = (($signed(_zz__31_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_24_inner_activation;
    end else begin
      io_macOut = _31_24_inner_macOut;
    end
  end

  assign _zz__31_24_inner_macOut = ($signed(_zz__zz__31_24_inner_macOut) + $signed(_zz__zz__31_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_24_inner_activation <= 8'h00;
      _31_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_24_inner_activation <= io_addInput;
      end else begin
        _31_24_inner_macOut <= _zz__31_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1015 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_23_inner_macOut;
  wire       [15:0]   _zz__zz__31_23_inner_macOut_1;
  wire       [15:0]   _zz__31_23_inner_macOut_1;
  wire       [15:0]   _zz__31_23_inner_macOut_2;
  reg        [7:0]    _31_23_inner_activation;
  reg        [7:0]    _31_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_23_inner_macOut;

  assign _zz__zz__31_23_inner_macOut = ($signed(io_mulInput) * $signed(_31_23_inner_activation));
  assign _zz__zz__31_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_23_inner_macOut)) ? 16'h007f : _zz__31_23_inner_macOut_2);
  assign _zz__31_23_inner_macOut_2 = (($signed(_zz__31_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_23_inner_activation;
    end else begin
      io_macOut = _31_23_inner_macOut;
    end
  end

  assign _zz__31_23_inner_macOut = ($signed(_zz__zz__31_23_inner_macOut) + $signed(_zz__zz__31_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_23_inner_activation <= 8'h00;
      _31_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_23_inner_activation <= io_addInput;
      end else begin
        _31_23_inner_macOut <= _zz__31_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1014 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_22_inner_macOut;
  wire       [15:0]   _zz__zz__31_22_inner_macOut_1;
  wire       [15:0]   _zz__31_22_inner_macOut_1;
  wire       [15:0]   _zz__31_22_inner_macOut_2;
  reg        [7:0]    _31_22_inner_activation;
  reg        [7:0]    _31_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_22_inner_macOut;

  assign _zz__zz__31_22_inner_macOut = ($signed(io_mulInput) * $signed(_31_22_inner_activation));
  assign _zz__zz__31_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_22_inner_macOut)) ? 16'h007f : _zz__31_22_inner_macOut_2);
  assign _zz__31_22_inner_macOut_2 = (($signed(_zz__31_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_22_inner_activation;
    end else begin
      io_macOut = _31_22_inner_macOut;
    end
  end

  assign _zz__31_22_inner_macOut = ($signed(_zz__zz__31_22_inner_macOut) + $signed(_zz__zz__31_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_22_inner_activation <= 8'h00;
      _31_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_22_inner_activation <= io_addInput;
      end else begin
        _31_22_inner_macOut <= _zz__31_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1013 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_21_inner_macOut;
  wire       [15:0]   _zz__zz__31_21_inner_macOut_1;
  wire       [15:0]   _zz__31_21_inner_macOut_1;
  wire       [15:0]   _zz__31_21_inner_macOut_2;
  reg        [7:0]    _31_21_inner_activation;
  reg        [7:0]    _31_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_21_inner_macOut;

  assign _zz__zz__31_21_inner_macOut = ($signed(io_mulInput) * $signed(_31_21_inner_activation));
  assign _zz__zz__31_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_21_inner_macOut)) ? 16'h007f : _zz__31_21_inner_macOut_2);
  assign _zz__31_21_inner_macOut_2 = (($signed(_zz__31_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_21_inner_activation;
    end else begin
      io_macOut = _31_21_inner_macOut;
    end
  end

  assign _zz__31_21_inner_macOut = ($signed(_zz__zz__31_21_inner_macOut) + $signed(_zz__zz__31_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_21_inner_activation <= 8'h00;
      _31_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_21_inner_activation <= io_addInput;
      end else begin
        _31_21_inner_macOut <= _zz__31_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1012 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_20_inner_macOut;
  wire       [15:0]   _zz__zz__31_20_inner_macOut_1;
  wire       [15:0]   _zz__31_20_inner_macOut_1;
  wire       [15:0]   _zz__31_20_inner_macOut_2;
  reg        [7:0]    _31_20_inner_activation;
  reg        [7:0]    _31_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_20_inner_macOut;

  assign _zz__zz__31_20_inner_macOut = ($signed(io_mulInput) * $signed(_31_20_inner_activation));
  assign _zz__zz__31_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_20_inner_macOut)) ? 16'h007f : _zz__31_20_inner_macOut_2);
  assign _zz__31_20_inner_macOut_2 = (($signed(_zz__31_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_20_inner_activation;
    end else begin
      io_macOut = _31_20_inner_macOut;
    end
  end

  assign _zz__31_20_inner_macOut = ($signed(_zz__zz__31_20_inner_macOut) + $signed(_zz__zz__31_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_20_inner_activation <= 8'h00;
      _31_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_20_inner_activation <= io_addInput;
      end else begin
        _31_20_inner_macOut <= _zz__31_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1011 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_19_inner_macOut;
  wire       [15:0]   _zz__zz__31_19_inner_macOut_1;
  wire       [15:0]   _zz__31_19_inner_macOut_1;
  wire       [15:0]   _zz__31_19_inner_macOut_2;
  reg        [7:0]    _31_19_inner_activation;
  reg        [7:0]    _31_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_19_inner_macOut;

  assign _zz__zz__31_19_inner_macOut = ($signed(io_mulInput) * $signed(_31_19_inner_activation));
  assign _zz__zz__31_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_19_inner_macOut)) ? 16'h007f : _zz__31_19_inner_macOut_2);
  assign _zz__31_19_inner_macOut_2 = (($signed(_zz__31_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_19_inner_activation;
    end else begin
      io_macOut = _31_19_inner_macOut;
    end
  end

  assign _zz__31_19_inner_macOut = ($signed(_zz__zz__31_19_inner_macOut) + $signed(_zz__zz__31_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_19_inner_activation <= 8'h00;
      _31_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_19_inner_activation <= io_addInput;
      end else begin
        _31_19_inner_macOut <= _zz__31_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1010 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_18_inner_macOut;
  wire       [15:0]   _zz__zz__31_18_inner_macOut_1;
  wire       [15:0]   _zz__31_18_inner_macOut_1;
  wire       [15:0]   _zz__31_18_inner_macOut_2;
  reg        [7:0]    _31_18_inner_activation;
  reg        [7:0]    _31_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_18_inner_macOut;

  assign _zz__zz__31_18_inner_macOut = ($signed(io_mulInput) * $signed(_31_18_inner_activation));
  assign _zz__zz__31_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_18_inner_macOut)) ? 16'h007f : _zz__31_18_inner_macOut_2);
  assign _zz__31_18_inner_macOut_2 = (($signed(_zz__31_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_18_inner_activation;
    end else begin
      io_macOut = _31_18_inner_macOut;
    end
  end

  assign _zz__31_18_inner_macOut = ($signed(_zz__zz__31_18_inner_macOut) + $signed(_zz__zz__31_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_18_inner_activation <= 8'h00;
      _31_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_18_inner_activation <= io_addInput;
      end else begin
        _31_18_inner_macOut <= _zz__31_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1009 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_17_inner_macOut;
  wire       [15:0]   _zz__zz__31_17_inner_macOut_1;
  wire       [15:0]   _zz__31_17_inner_macOut_1;
  wire       [15:0]   _zz__31_17_inner_macOut_2;
  reg        [7:0]    _31_17_inner_activation;
  reg        [7:0]    _31_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_17_inner_macOut;

  assign _zz__zz__31_17_inner_macOut = ($signed(io_mulInput) * $signed(_31_17_inner_activation));
  assign _zz__zz__31_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_17_inner_macOut)) ? 16'h007f : _zz__31_17_inner_macOut_2);
  assign _zz__31_17_inner_macOut_2 = (($signed(_zz__31_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_17_inner_activation;
    end else begin
      io_macOut = _31_17_inner_macOut;
    end
  end

  assign _zz__31_17_inner_macOut = ($signed(_zz__zz__31_17_inner_macOut) + $signed(_zz__zz__31_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_17_inner_activation <= 8'h00;
      _31_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_17_inner_activation <= io_addInput;
      end else begin
        _31_17_inner_macOut <= _zz__31_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1008 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_16_inner_macOut;
  wire       [15:0]   _zz__zz__31_16_inner_macOut_1;
  wire       [15:0]   _zz__31_16_inner_macOut_1;
  wire       [15:0]   _zz__31_16_inner_macOut_2;
  reg        [7:0]    _31_16_inner_activation;
  reg        [7:0]    _31_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_16_inner_macOut;

  assign _zz__zz__31_16_inner_macOut = ($signed(io_mulInput) * $signed(_31_16_inner_activation));
  assign _zz__zz__31_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_16_inner_macOut)) ? 16'h007f : _zz__31_16_inner_macOut_2);
  assign _zz__31_16_inner_macOut_2 = (($signed(_zz__31_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_16_inner_activation;
    end else begin
      io_macOut = _31_16_inner_macOut;
    end
  end

  assign _zz__31_16_inner_macOut = ($signed(_zz__zz__31_16_inner_macOut) + $signed(_zz__zz__31_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_16_inner_activation <= 8'h00;
      _31_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_16_inner_activation <= io_addInput;
      end else begin
        _31_16_inner_macOut <= _zz__31_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1007 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_15_inner_macOut;
  wire       [15:0]   _zz__zz__31_15_inner_macOut_1;
  wire       [15:0]   _zz__31_15_inner_macOut_1;
  wire       [15:0]   _zz__31_15_inner_macOut_2;
  reg        [7:0]    _31_15_inner_activation;
  reg        [7:0]    _31_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_15_inner_macOut;

  assign _zz__zz__31_15_inner_macOut = ($signed(io_mulInput) * $signed(_31_15_inner_activation));
  assign _zz__zz__31_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_15_inner_macOut)) ? 16'h007f : _zz__31_15_inner_macOut_2);
  assign _zz__31_15_inner_macOut_2 = (($signed(_zz__31_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_15_inner_activation;
    end else begin
      io_macOut = _31_15_inner_macOut;
    end
  end

  assign _zz__31_15_inner_macOut = ($signed(_zz__zz__31_15_inner_macOut) + $signed(_zz__zz__31_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_15_inner_activation <= 8'h00;
      _31_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_15_inner_activation <= io_addInput;
      end else begin
        _31_15_inner_macOut <= _zz__31_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1006 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_14_inner_macOut;
  wire       [15:0]   _zz__zz__31_14_inner_macOut_1;
  wire       [15:0]   _zz__31_14_inner_macOut_1;
  wire       [15:0]   _zz__31_14_inner_macOut_2;
  reg        [7:0]    _31_14_inner_activation;
  reg        [7:0]    _31_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_14_inner_macOut;

  assign _zz__zz__31_14_inner_macOut = ($signed(io_mulInput) * $signed(_31_14_inner_activation));
  assign _zz__zz__31_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_14_inner_macOut)) ? 16'h007f : _zz__31_14_inner_macOut_2);
  assign _zz__31_14_inner_macOut_2 = (($signed(_zz__31_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_14_inner_activation;
    end else begin
      io_macOut = _31_14_inner_macOut;
    end
  end

  assign _zz__31_14_inner_macOut = ($signed(_zz__zz__31_14_inner_macOut) + $signed(_zz__zz__31_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_14_inner_activation <= 8'h00;
      _31_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_14_inner_activation <= io_addInput;
      end else begin
        _31_14_inner_macOut <= _zz__31_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1005 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_13_inner_macOut;
  wire       [15:0]   _zz__zz__31_13_inner_macOut_1;
  wire       [15:0]   _zz__31_13_inner_macOut_1;
  wire       [15:0]   _zz__31_13_inner_macOut_2;
  reg        [7:0]    _31_13_inner_activation;
  reg        [7:0]    _31_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_13_inner_macOut;

  assign _zz__zz__31_13_inner_macOut = ($signed(io_mulInput) * $signed(_31_13_inner_activation));
  assign _zz__zz__31_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_13_inner_macOut)) ? 16'h007f : _zz__31_13_inner_macOut_2);
  assign _zz__31_13_inner_macOut_2 = (($signed(_zz__31_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_13_inner_activation;
    end else begin
      io_macOut = _31_13_inner_macOut;
    end
  end

  assign _zz__31_13_inner_macOut = ($signed(_zz__zz__31_13_inner_macOut) + $signed(_zz__zz__31_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_13_inner_activation <= 8'h00;
      _31_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_13_inner_activation <= io_addInput;
      end else begin
        _31_13_inner_macOut <= _zz__31_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1004 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_12_inner_macOut;
  wire       [15:0]   _zz__zz__31_12_inner_macOut_1;
  wire       [15:0]   _zz__31_12_inner_macOut_1;
  wire       [15:0]   _zz__31_12_inner_macOut_2;
  reg        [7:0]    _31_12_inner_activation;
  reg        [7:0]    _31_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_12_inner_macOut;

  assign _zz__zz__31_12_inner_macOut = ($signed(io_mulInput) * $signed(_31_12_inner_activation));
  assign _zz__zz__31_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_12_inner_macOut)) ? 16'h007f : _zz__31_12_inner_macOut_2);
  assign _zz__31_12_inner_macOut_2 = (($signed(_zz__31_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_12_inner_activation;
    end else begin
      io_macOut = _31_12_inner_macOut;
    end
  end

  assign _zz__31_12_inner_macOut = ($signed(_zz__zz__31_12_inner_macOut) + $signed(_zz__zz__31_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_12_inner_activation <= 8'h00;
      _31_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_12_inner_activation <= io_addInput;
      end else begin
        _31_12_inner_macOut <= _zz__31_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1003 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_11_inner_macOut;
  wire       [15:0]   _zz__zz__31_11_inner_macOut_1;
  wire       [15:0]   _zz__31_11_inner_macOut_1;
  wire       [15:0]   _zz__31_11_inner_macOut_2;
  reg        [7:0]    _31_11_inner_activation;
  reg        [7:0]    _31_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_11_inner_macOut;

  assign _zz__zz__31_11_inner_macOut = ($signed(io_mulInput) * $signed(_31_11_inner_activation));
  assign _zz__zz__31_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_11_inner_macOut)) ? 16'h007f : _zz__31_11_inner_macOut_2);
  assign _zz__31_11_inner_macOut_2 = (($signed(_zz__31_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_11_inner_activation;
    end else begin
      io_macOut = _31_11_inner_macOut;
    end
  end

  assign _zz__31_11_inner_macOut = ($signed(_zz__zz__31_11_inner_macOut) + $signed(_zz__zz__31_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_11_inner_activation <= 8'h00;
      _31_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_11_inner_activation <= io_addInput;
      end else begin
        _31_11_inner_macOut <= _zz__31_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1002 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_10_inner_macOut;
  wire       [15:0]   _zz__zz__31_10_inner_macOut_1;
  wire       [15:0]   _zz__31_10_inner_macOut_1;
  wire       [15:0]   _zz__31_10_inner_macOut_2;
  reg        [7:0]    _31_10_inner_activation;
  reg        [7:0]    _31_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_10_inner_macOut;

  assign _zz__zz__31_10_inner_macOut = ($signed(io_mulInput) * $signed(_31_10_inner_activation));
  assign _zz__zz__31_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_10_inner_macOut)) ? 16'h007f : _zz__31_10_inner_macOut_2);
  assign _zz__31_10_inner_macOut_2 = (($signed(_zz__31_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_10_inner_activation;
    end else begin
      io_macOut = _31_10_inner_macOut;
    end
  end

  assign _zz__31_10_inner_macOut = ($signed(_zz__zz__31_10_inner_macOut) + $signed(_zz__zz__31_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_10_inner_activation <= 8'h00;
      _31_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_10_inner_activation <= io_addInput;
      end else begin
        _31_10_inner_macOut <= _zz__31_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1001 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_9_inner_macOut;
  wire       [15:0]   _zz__zz__31_9_inner_macOut_1;
  wire       [15:0]   _zz__31_9_inner_macOut_1;
  wire       [15:0]   _zz__31_9_inner_macOut_2;
  reg        [7:0]    _31_9_inner_activation;
  reg        [7:0]    _31_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_9_inner_macOut;

  assign _zz__zz__31_9_inner_macOut = ($signed(io_mulInput) * $signed(_31_9_inner_activation));
  assign _zz__zz__31_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_9_inner_macOut)) ? 16'h007f : _zz__31_9_inner_macOut_2);
  assign _zz__31_9_inner_macOut_2 = (($signed(_zz__31_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_9_inner_activation;
    end else begin
      io_macOut = _31_9_inner_macOut;
    end
  end

  assign _zz__31_9_inner_macOut = ($signed(_zz__zz__31_9_inner_macOut) + $signed(_zz__zz__31_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_9_inner_activation <= 8'h00;
      _31_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_9_inner_activation <= io_addInput;
      end else begin
        _31_9_inner_macOut <= _zz__31_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1000 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_8_inner_macOut;
  wire       [15:0]   _zz__zz__31_8_inner_macOut_1;
  wire       [15:0]   _zz__31_8_inner_macOut_1;
  wire       [15:0]   _zz__31_8_inner_macOut_2;
  reg        [7:0]    _31_8_inner_activation;
  reg        [7:0]    _31_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_8_inner_macOut;

  assign _zz__zz__31_8_inner_macOut = ($signed(io_mulInput) * $signed(_31_8_inner_activation));
  assign _zz__zz__31_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_8_inner_macOut)) ? 16'h007f : _zz__31_8_inner_macOut_2);
  assign _zz__31_8_inner_macOut_2 = (($signed(_zz__31_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_8_inner_activation;
    end else begin
      io_macOut = _31_8_inner_macOut;
    end
  end

  assign _zz__31_8_inner_macOut = ($signed(_zz__zz__31_8_inner_macOut) + $signed(_zz__zz__31_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_8_inner_activation <= 8'h00;
      _31_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_8_inner_activation <= io_addInput;
      end else begin
        _31_8_inner_macOut <= _zz__31_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_999 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_7_inner_macOut;
  wire       [15:0]   _zz__zz__31_7_inner_macOut_1;
  wire       [15:0]   _zz__31_7_inner_macOut_1;
  wire       [15:0]   _zz__31_7_inner_macOut_2;
  reg        [7:0]    _31_7_inner_activation;
  reg        [7:0]    _31_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_7_inner_macOut;

  assign _zz__zz__31_7_inner_macOut = ($signed(io_mulInput) * $signed(_31_7_inner_activation));
  assign _zz__zz__31_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_7_inner_macOut)) ? 16'h007f : _zz__31_7_inner_macOut_2);
  assign _zz__31_7_inner_macOut_2 = (($signed(_zz__31_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_7_inner_activation;
    end else begin
      io_macOut = _31_7_inner_macOut;
    end
  end

  assign _zz__31_7_inner_macOut = ($signed(_zz__zz__31_7_inner_macOut) + $signed(_zz__zz__31_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_7_inner_activation <= 8'h00;
      _31_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_7_inner_activation <= io_addInput;
      end else begin
        _31_7_inner_macOut <= _zz__31_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_998 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_6_inner_macOut;
  wire       [15:0]   _zz__zz__31_6_inner_macOut_1;
  wire       [15:0]   _zz__31_6_inner_macOut_1;
  wire       [15:0]   _zz__31_6_inner_macOut_2;
  reg        [7:0]    _31_6_inner_activation;
  reg        [7:0]    _31_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_6_inner_macOut;

  assign _zz__zz__31_6_inner_macOut = ($signed(io_mulInput) * $signed(_31_6_inner_activation));
  assign _zz__zz__31_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_6_inner_macOut)) ? 16'h007f : _zz__31_6_inner_macOut_2);
  assign _zz__31_6_inner_macOut_2 = (($signed(_zz__31_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_6_inner_activation;
    end else begin
      io_macOut = _31_6_inner_macOut;
    end
  end

  assign _zz__31_6_inner_macOut = ($signed(_zz__zz__31_6_inner_macOut) + $signed(_zz__zz__31_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_6_inner_activation <= 8'h00;
      _31_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_6_inner_activation <= io_addInput;
      end else begin
        _31_6_inner_macOut <= _zz__31_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_997 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_5_inner_macOut;
  wire       [15:0]   _zz__zz__31_5_inner_macOut_1;
  wire       [15:0]   _zz__31_5_inner_macOut_1;
  wire       [15:0]   _zz__31_5_inner_macOut_2;
  reg        [7:0]    _31_5_inner_activation;
  reg        [7:0]    _31_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_5_inner_macOut;

  assign _zz__zz__31_5_inner_macOut = ($signed(io_mulInput) * $signed(_31_5_inner_activation));
  assign _zz__zz__31_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_5_inner_macOut)) ? 16'h007f : _zz__31_5_inner_macOut_2);
  assign _zz__31_5_inner_macOut_2 = (($signed(_zz__31_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_5_inner_activation;
    end else begin
      io_macOut = _31_5_inner_macOut;
    end
  end

  assign _zz__31_5_inner_macOut = ($signed(_zz__zz__31_5_inner_macOut) + $signed(_zz__zz__31_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_5_inner_activation <= 8'h00;
      _31_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_5_inner_activation <= io_addInput;
      end else begin
        _31_5_inner_macOut <= _zz__31_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_996 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_4_inner_macOut;
  wire       [15:0]   _zz__zz__31_4_inner_macOut_1;
  wire       [15:0]   _zz__31_4_inner_macOut_1;
  wire       [15:0]   _zz__31_4_inner_macOut_2;
  reg        [7:0]    _31_4_inner_activation;
  reg        [7:0]    _31_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_4_inner_macOut;

  assign _zz__zz__31_4_inner_macOut = ($signed(io_mulInput) * $signed(_31_4_inner_activation));
  assign _zz__zz__31_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_4_inner_macOut)) ? 16'h007f : _zz__31_4_inner_macOut_2);
  assign _zz__31_4_inner_macOut_2 = (($signed(_zz__31_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_4_inner_activation;
    end else begin
      io_macOut = _31_4_inner_macOut;
    end
  end

  assign _zz__31_4_inner_macOut = ($signed(_zz__zz__31_4_inner_macOut) + $signed(_zz__zz__31_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_4_inner_activation <= 8'h00;
      _31_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_4_inner_activation <= io_addInput;
      end else begin
        _31_4_inner_macOut <= _zz__31_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_995 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_3_inner_macOut;
  wire       [15:0]   _zz__zz__31_3_inner_macOut_1;
  wire       [15:0]   _zz__31_3_inner_macOut_1;
  wire       [15:0]   _zz__31_3_inner_macOut_2;
  reg        [7:0]    _31_3_inner_activation;
  reg        [7:0]    _31_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_3_inner_macOut;

  assign _zz__zz__31_3_inner_macOut = ($signed(io_mulInput) * $signed(_31_3_inner_activation));
  assign _zz__zz__31_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_3_inner_macOut)) ? 16'h007f : _zz__31_3_inner_macOut_2);
  assign _zz__31_3_inner_macOut_2 = (($signed(_zz__31_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_3_inner_activation;
    end else begin
      io_macOut = _31_3_inner_macOut;
    end
  end

  assign _zz__31_3_inner_macOut = ($signed(_zz__zz__31_3_inner_macOut) + $signed(_zz__zz__31_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_3_inner_activation <= 8'h00;
      _31_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_3_inner_activation <= io_addInput;
      end else begin
        _31_3_inner_macOut <= _zz__31_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_994 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_2_inner_macOut;
  wire       [15:0]   _zz__zz__31_2_inner_macOut_1;
  wire       [15:0]   _zz__31_2_inner_macOut_1;
  wire       [15:0]   _zz__31_2_inner_macOut_2;
  reg        [7:0]    _31_2_inner_activation;
  reg        [7:0]    _31_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_2_inner_macOut;

  assign _zz__zz__31_2_inner_macOut = ($signed(io_mulInput) * $signed(_31_2_inner_activation));
  assign _zz__zz__31_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_2_inner_macOut)) ? 16'h007f : _zz__31_2_inner_macOut_2);
  assign _zz__31_2_inner_macOut_2 = (($signed(_zz__31_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_2_inner_activation;
    end else begin
      io_macOut = _31_2_inner_macOut;
    end
  end

  assign _zz__31_2_inner_macOut = ($signed(_zz__zz__31_2_inner_macOut) + $signed(_zz__zz__31_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_2_inner_activation <= 8'h00;
      _31_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_2_inner_activation <= io_addInput;
      end else begin
        _31_2_inner_macOut <= _zz__31_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_993 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_1_inner_macOut;
  wire       [15:0]   _zz__zz__31_1_inner_macOut_1;
  wire       [15:0]   _zz__31_1_inner_macOut_1;
  wire       [15:0]   _zz__31_1_inner_macOut_2;
  reg        [7:0]    _31_1_inner_activation;
  reg        [7:0]    _31_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_1_inner_macOut;

  assign _zz__zz__31_1_inner_macOut = ($signed(io_mulInput) * $signed(_31_1_inner_activation));
  assign _zz__zz__31_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_1_inner_macOut)) ? 16'h007f : _zz__31_1_inner_macOut_2);
  assign _zz__31_1_inner_macOut_2 = (($signed(_zz__31_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_1_inner_activation;
    end else begin
      io_macOut = _31_1_inner_macOut;
    end
  end

  assign _zz__31_1_inner_macOut = ($signed(_zz__zz__31_1_inner_macOut) + $signed(_zz__zz__31_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_1_inner_activation <= 8'h00;
      _31_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_1_inner_activation <= io_addInput;
      end else begin
        _31_1_inner_macOut <= _zz__31_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_992 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__31_0_inner_macOut;
  wire       [15:0]   _zz__zz__31_0_inner_macOut_1;
  wire       [15:0]   _zz__31_0_inner_macOut_1;
  wire       [15:0]   _zz__31_0_inner_macOut_2;
  reg        [7:0]    _31_0_inner_activation;
  reg        [7:0]    _31_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__31_0_inner_macOut;

  assign _zz__zz__31_0_inner_macOut = ($signed(io_mulInput) * $signed(_31_0_inner_activation));
  assign _zz__zz__31_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__31_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__31_0_inner_macOut)) ? 16'h007f : _zz__31_0_inner_macOut_2);
  assign _zz__31_0_inner_macOut_2 = (($signed(_zz__31_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__31_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _31_0_inner_activation;
    end else begin
      io_macOut = _31_0_inner_macOut;
    end
  end

  assign _zz__31_0_inner_macOut = ($signed(_zz__zz__31_0_inner_macOut) + $signed(_zz__zz__31_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _31_0_inner_activation <= 8'h00;
      _31_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _31_0_inner_activation <= io_addInput;
      end else begin
        _31_0_inner_macOut <= _zz__31_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_991 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_31_inner_macOut;
  wire       [15:0]   _zz__zz__30_31_inner_macOut_1;
  wire       [15:0]   _zz__30_31_inner_macOut_1;
  wire       [15:0]   _zz__30_31_inner_macOut_2;
  reg        [7:0]    _30_31_inner_activation;
  reg        [7:0]    _30_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_31_inner_macOut;

  assign _zz__zz__30_31_inner_macOut = ($signed(io_mulInput) * $signed(_30_31_inner_activation));
  assign _zz__zz__30_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_31_inner_macOut)) ? 16'h007f : _zz__30_31_inner_macOut_2);
  assign _zz__30_31_inner_macOut_2 = (($signed(_zz__30_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_31_inner_activation;
    end else begin
      io_macOut = _30_31_inner_macOut;
    end
  end

  assign _zz__30_31_inner_macOut = ($signed(_zz__zz__30_31_inner_macOut) + $signed(_zz__zz__30_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_31_inner_activation <= 8'h00;
      _30_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_31_inner_activation <= io_addInput;
      end else begin
        _30_31_inner_macOut <= _zz__30_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_990 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_30_inner_macOut;
  wire       [15:0]   _zz__zz__30_30_inner_macOut_1;
  wire       [15:0]   _zz__30_30_inner_macOut_1;
  wire       [15:0]   _zz__30_30_inner_macOut_2;
  reg        [7:0]    _30_30_inner_activation;
  reg        [7:0]    _30_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_30_inner_macOut;

  assign _zz__zz__30_30_inner_macOut = ($signed(io_mulInput) * $signed(_30_30_inner_activation));
  assign _zz__zz__30_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_30_inner_macOut)) ? 16'h007f : _zz__30_30_inner_macOut_2);
  assign _zz__30_30_inner_macOut_2 = (($signed(_zz__30_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_30_inner_activation;
    end else begin
      io_macOut = _30_30_inner_macOut;
    end
  end

  assign _zz__30_30_inner_macOut = ($signed(_zz__zz__30_30_inner_macOut) + $signed(_zz__zz__30_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_30_inner_activation <= 8'h00;
      _30_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_30_inner_activation <= io_addInput;
      end else begin
        _30_30_inner_macOut <= _zz__30_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_989 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_29_inner_macOut;
  wire       [15:0]   _zz__zz__30_29_inner_macOut_1;
  wire       [15:0]   _zz__30_29_inner_macOut_1;
  wire       [15:0]   _zz__30_29_inner_macOut_2;
  reg        [7:0]    _30_29_inner_activation;
  reg        [7:0]    _30_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_29_inner_macOut;

  assign _zz__zz__30_29_inner_macOut = ($signed(io_mulInput) * $signed(_30_29_inner_activation));
  assign _zz__zz__30_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_29_inner_macOut)) ? 16'h007f : _zz__30_29_inner_macOut_2);
  assign _zz__30_29_inner_macOut_2 = (($signed(_zz__30_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_29_inner_activation;
    end else begin
      io_macOut = _30_29_inner_macOut;
    end
  end

  assign _zz__30_29_inner_macOut = ($signed(_zz__zz__30_29_inner_macOut) + $signed(_zz__zz__30_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_29_inner_activation <= 8'h00;
      _30_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_29_inner_activation <= io_addInput;
      end else begin
        _30_29_inner_macOut <= _zz__30_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_988 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_28_inner_macOut;
  wire       [15:0]   _zz__zz__30_28_inner_macOut_1;
  wire       [15:0]   _zz__30_28_inner_macOut_1;
  wire       [15:0]   _zz__30_28_inner_macOut_2;
  reg        [7:0]    _30_28_inner_activation;
  reg        [7:0]    _30_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_28_inner_macOut;

  assign _zz__zz__30_28_inner_macOut = ($signed(io_mulInput) * $signed(_30_28_inner_activation));
  assign _zz__zz__30_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_28_inner_macOut)) ? 16'h007f : _zz__30_28_inner_macOut_2);
  assign _zz__30_28_inner_macOut_2 = (($signed(_zz__30_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_28_inner_activation;
    end else begin
      io_macOut = _30_28_inner_macOut;
    end
  end

  assign _zz__30_28_inner_macOut = ($signed(_zz__zz__30_28_inner_macOut) + $signed(_zz__zz__30_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_28_inner_activation <= 8'h00;
      _30_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_28_inner_activation <= io_addInput;
      end else begin
        _30_28_inner_macOut <= _zz__30_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_987 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_27_inner_macOut;
  wire       [15:0]   _zz__zz__30_27_inner_macOut_1;
  wire       [15:0]   _zz__30_27_inner_macOut_1;
  wire       [15:0]   _zz__30_27_inner_macOut_2;
  reg        [7:0]    _30_27_inner_activation;
  reg        [7:0]    _30_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_27_inner_macOut;

  assign _zz__zz__30_27_inner_macOut = ($signed(io_mulInput) * $signed(_30_27_inner_activation));
  assign _zz__zz__30_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_27_inner_macOut)) ? 16'h007f : _zz__30_27_inner_macOut_2);
  assign _zz__30_27_inner_macOut_2 = (($signed(_zz__30_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_27_inner_activation;
    end else begin
      io_macOut = _30_27_inner_macOut;
    end
  end

  assign _zz__30_27_inner_macOut = ($signed(_zz__zz__30_27_inner_macOut) + $signed(_zz__zz__30_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_27_inner_activation <= 8'h00;
      _30_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_27_inner_activation <= io_addInput;
      end else begin
        _30_27_inner_macOut <= _zz__30_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_986 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_26_inner_macOut;
  wire       [15:0]   _zz__zz__30_26_inner_macOut_1;
  wire       [15:0]   _zz__30_26_inner_macOut_1;
  wire       [15:0]   _zz__30_26_inner_macOut_2;
  reg        [7:0]    _30_26_inner_activation;
  reg        [7:0]    _30_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_26_inner_macOut;

  assign _zz__zz__30_26_inner_macOut = ($signed(io_mulInput) * $signed(_30_26_inner_activation));
  assign _zz__zz__30_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_26_inner_macOut)) ? 16'h007f : _zz__30_26_inner_macOut_2);
  assign _zz__30_26_inner_macOut_2 = (($signed(_zz__30_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_26_inner_activation;
    end else begin
      io_macOut = _30_26_inner_macOut;
    end
  end

  assign _zz__30_26_inner_macOut = ($signed(_zz__zz__30_26_inner_macOut) + $signed(_zz__zz__30_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_26_inner_activation <= 8'h00;
      _30_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_26_inner_activation <= io_addInput;
      end else begin
        _30_26_inner_macOut <= _zz__30_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_985 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_25_inner_macOut;
  wire       [15:0]   _zz__zz__30_25_inner_macOut_1;
  wire       [15:0]   _zz__30_25_inner_macOut_1;
  wire       [15:0]   _zz__30_25_inner_macOut_2;
  reg        [7:0]    _30_25_inner_activation;
  reg        [7:0]    _30_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_25_inner_macOut;

  assign _zz__zz__30_25_inner_macOut = ($signed(io_mulInput) * $signed(_30_25_inner_activation));
  assign _zz__zz__30_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_25_inner_macOut)) ? 16'h007f : _zz__30_25_inner_macOut_2);
  assign _zz__30_25_inner_macOut_2 = (($signed(_zz__30_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_25_inner_activation;
    end else begin
      io_macOut = _30_25_inner_macOut;
    end
  end

  assign _zz__30_25_inner_macOut = ($signed(_zz__zz__30_25_inner_macOut) + $signed(_zz__zz__30_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_25_inner_activation <= 8'h00;
      _30_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_25_inner_activation <= io_addInput;
      end else begin
        _30_25_inner_macOut <= _zz__30_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_984 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_24_inner_macOut;
  wire       [15:0]   _zz__zz__30_24_inner_macOut_1;
  wire       [15:0]   _zz__30_24_inner_macOut_1;
  wire       [15:0]   _zz__30_24_inner_macOut_2;
  reg        [7:0]    _30_24_inner_activation;
  reg        [7:0]    _30_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_24_inner_macOut;

  assign _zz__zz__30_24_inner_macOut = ($signed(io_mulInput) * $signed(_30_24_inner_activation));
  assign _zz__zz__30_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_24_inner_macOut)) ? 16'h007f : _zz__30_24_inner_macOut_2);
  assign _zz__30_24_inner_macOut_2 = (($signed(_zz__30_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_24_inner_activation;
    end else begin
      io_macOut = _30_24_inner_macOut;
    end
  end

  assign _zz__30_24_inner_macOut = ($signed(_zz__zz__30_24_inner_macOut) + $signed(_zz__zz__30_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_24_inner_activation <= 8'h00;
      _30_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_24_inner_activation <= io_addInput;
      end else begin
        _30_24_inner_macOut <= _zz__30_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_983 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_23_inner_macOut;
  wire       [15:0]   _zz__zz__30_23_inner_macOut_1;
  wire       [15:0]   _zz__30_23_inner_macOut_1;
  wire       [15:0]   _zz__30_23_inner_macOut_2;
  reg        [7:0]    _30_23_inner_activation;
  reg        [7:0]    _30_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_23_inner_macOut;

  assign _zz__zz__30_23_inner_macOut = ($signed(io_mulInput) * $signed(_30_23_inner_activation));
  assign _zz__zz__30_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_23_inner_macOut)) ? 16'h007f : _zz__30_23_inner_macOut_2);
  assign _zz__30_23_inner_macOut_2 = (($signed(_zz__30_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_23_inner_activation;
    end else begin
      io_macOut = _30_23_inner_macOut;
    end
  end

  assign _zz__30_23_inner_macOut = ($signed(_zz__zz__30_23_inner_macOut) + $signed(_zz__zz__30_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_23_inner_activation <= 8'h00;
      _30_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_23_inner_activation <= io_addInput;
      end else begin
        _30_23_inner_macOut <= _zz__30_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_982 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_22_inner_macOut;
  wire       [15:0]   _zz__zz__30_22_inner_macOut_1;
  wire       [15:0]   _zz__30_22_inner_macOut_1;
  wire       [15:0]   _zz__30_22_inner_macOut_2;
  reg        [7:0]    _30_22_inner_activation;
  reg        [7:0]    _30_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_22_inner_macOut;

  assign _zz__zz__30_22_inner_macOut = ($signed(io_mulInput) * $signed(_30_22_inner_activation));
  assign _zz__zz__30_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_22_inner_macOut)) ? 16'h007f : _zz__30_22_inner_macOut_2);
  assign _zz__30_22_inner_macOut_2 = (($signed(_zz__30_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_22_inner_activation;
    end else begin
      io_macOut = _30_22_inner_macOut;
    end
  end

  assign _zz__30_22_inner_macOut = ($signed(_zz__zz__30_22_inner_macOut) + $signed(_zz__zz__30_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_22_inner_activation <= 8'h00;
      _30_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_22_inner_activation <= io_addInput;
      end else begin
        _30_22_inner_macOut <= _zz__30_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_981 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_21_inner_macOut;
  wire       [15:0]   _zz__zz__30_21_inner_macOut_1;
  wire       [15:0]   _zz__30_21_inner_macOut_1;
  wire       [15:0]   _zz__30_21_inner_macOut_2;
  reg        [7:0]    _30_21_inner_activation;
  reg        [7:0]    _30_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_21_inner_macOut;

  assign _zz__zz__30_21_inner_macOut = ($signed(io_mulInput) * $signed(_30_21_inner_activation));
  assign _zz__zz__30_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_21_inner_macOut)) ? 16'h007f : _zz__30_21_inner_macOut_2);
  assign _zz__30_21_inner_macOut_2 = (($signed(_zz__30_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_21_inner_activation;
    end else begin
      io_macOut = _30_21_inner_macOut;
    end
  end

  assign _zz__30_21_inner_macOut = ($signed(_zz__zz__30_21_inner_macOut) + $signed(_zz__zz__30_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_21_inner_activation <= 8'h00;
      _30_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_21_inner_activation <= io_addInput;
      end else begin
        _30_21_inner_macOut <= _zz__30_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_980 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_20_inner_macOut;
  wire       [15:0]   _zz__zz__30_20_inner_macOut_1;
  wire       [15:0]   _zz__30_20_inner_macOut_1;
  wire       [15:0]   _zz__30_20_inner_macOut_2;
  reg        [7:0]    _30_20_inner_activation;
  reg        [7:0]    _30_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_20_inner_macOut;

  assign _zz__zz__30_20_inner_macOut = ($signed(io_mulInput) * $signed(_30_20_inner_activation));
  assign _zz__zz__30_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_20_inner_macOut)) ? 16'h007f : _zz__30_20_inner_macOut_2);
  assign _zz__30_20_inner_macOut_2 = (($signed(_zz__30_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_20_inner_activation;
    end else begin
      io_macOut = _30_20_inner_macOut;
    end
  end

  assign _zz__30_20_inner_macOut = ($signed(_zz__zz__30_20_inner_macOut) + $signed(_zz__zz__30_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_20_inner_activation <= 8'h00;
      _30_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_20_inner_activation <= io_addInput;
      end else begin
        _30_20_inner_macOut <= _zz__30_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_979 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_19_inner_macOut;
  wire       [15:0]   _zz__zz__30_19_inner_macOut_1;
  wire       [15:0]   _zz__30_19_inner_macOut_1;
  wire       [15:0]   _zz__30_19_inner_macOut_2;
  reg        [7:0]    _30_19_inner_activation;
  reg        [7:0]    _30_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_19_inner_macOut;

  assign _zz__zz__30_19_inner_macOut = ($signed(io_mulInput) * $signed(_30_19_inner_activation));
  assign _zz__zz__30_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_19_inner_macOut)) ? 16'h007f : _zz__30_19_inner_macOut_2);
  assign _zz__30_19_inner_macOut_2 = (($signed(_zz__30_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_19_inner_activation;
    end else begin
      io_macOut = _30_19_inner_macOut;
    end
  end

  assign _zz__30_19_inner_macOut = ($signed(_zz__zz__30_19_inner_macOut) + $signed(_zz__zz__30_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_19_inner_activation <= 8'h00;
      _30_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_19_inner_activation <= io_addInput;
      end else begin
        _30_19_inner_macOut <= _zz__30_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_978 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_18_inner_macOut;
  wire       [15:0]   _zz__zz__30_18_inner_macOut_1;
  wire       [15:0]   _zz__30_18_inner_macOut_1;
  wire       [15:0]   _zz__30_18_inner_macOut_2;
  reg        [7:0]    _30_18_inner_activation;
  reg        [7:0]    _30_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_18_inner_macOut;

  assign _zz__zz__30_18_inner_macOut = ($signed(io_mulInput) * $signed(_30_18_inner_activation));
  assign _zz__zz__30_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_18_inner_macOut)) ? 16'h007f : _zz__30_18_inner_macOut_2);
  assign _zz__30_18_inner_macOut_2 = (($signed(_zz__30_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_18_inner_activation;
    end else begin
      io_macOut = _30_18_inner_macOut;
    end
  end

  assign _zz__30_18_inner_macOut = ($signed(_zz__zz__30_18_inner_macOut) + $signed(_zz__zz__30_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_18_inner_activation <= 8'h00;
      _30_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_18_inner_activation <= io_addInput;
      end else begin
        _30_18_inner_macOut <= _zz__30_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_977 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_17_inner_macOut;
  wire       [15:0]   _zz__zz__30_17_inner_macOut_1;
  wire       [15:0]   _zz__30_17_inner_macOut_1;
  wire       [15:0]   _zz__30_17_inner_macOut_2;
  reg        [7:0]    _30_17_inner_activation;
  reg        [7:0]    _30_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_17_inner_macOut;

  assign _zz__zz__30_17_inner_macOut = ($signed(io_mulInput) * $signed(_30_17_inner_activation));
  assign _zz__zz__30_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_17_inner_macOut)) ? 16'h007f : _zz__30_17_inner_macOut_2);
  assign _zz__30_17_inner_macOut_2 = (($signed(_zz__30_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_17_inner_activation;
    end else begin
      io_macOut = _30_17_inner_macOut;
    end
  end

  assign _zz__30_17_inner_macOut = ($signed(_zz__zz__30_17_inner_macOut) + $signed(_zz__zz__30_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_17_inner_activation <= 8'h00;
      _30_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_17_inner_activation <= io_addInput;
      end else begin
        _30_17_inner_macOut <= _zz__30_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_976 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_16_inner_macOut;
  wire       [15:0]   _zz__zz__30_16_inner_macOut_1;
  wire       [15:0]   _zz__30_16_inner_macOut_1;
  wire       [15:0]   _zz__30_16_inner_macOut_2;
  reg        [7:0]    _30_16_inner_activation;
  reg        [7:0]    _30_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_16_inner_macOut;

  assign _zz__zz__30_16_inner_macOut = ($signed(io_mulInput) * $signed(_30_16_inner_activation));
  assign _zz__zz__30_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_16_inner_macOut)) ? 16'h007f : _zz__30_16_inner_macOut_2);
  assign _zz__30_16_inner_macOut_2 = (($signed(_zz__30_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_16_inner_activation;
    end else begin
      io_macOut = _30_16_inner_macOut;
    end
  end

  assign _zz__30_16_inner_macOut = ($signed(_zz__zz__30_16_inner_macOut) + $signed(_zz__zz__30_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_16_inner_activation <= 8'h00;
      _30_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_16_inner_activation <= io_addInput;
      end else begin
        _30_16_inner_macOut <= _zz__30_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_975 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_15_inner_macOut;
  wire       [15:0]   _zz__zz__30_15_inner_macOut_1;
  wire       [15:0]   _zz__30_15_inner_macOut_1;
  wire       [15:0]   _zz__30_15_inner_macOut_2;
  reg        [7:0]    _30_15_inner_activation;
  reg        [7:0]    _30_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_15_inner_macOut;

  assign _zz__zz__30_15_inner_macOut = ($signed(io_mulInput) * $signed(_30_15_inner_activation));
  assign _zz__zz__30_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_15_inner_macOut)) ? 16'h007f : _zz__30_15_inner_macOut_2);
  assign _zz__30_15_inner_macOut_2 = (($signed(_zz__30_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_15_inner_activation;
    end else begin
      io_macOut = _30_15_inner_macOut;
    end
  end

  assign _zz__30_15_inner_macOut = ($signed(_zz__zz__30_15_inner_macOut) + $signed(_zz__zz__30_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_15_inner_activation <= 8'h00;
      _30_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_15_inner_activation <= io_addInput;
      end else begin
        _30_15_inner_macOut <= _zz__30_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_974 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_14_inner_macOut;
  wire       [15:0]   _zz__zz__30_14_inner_macOut_1;
  wire       [15:0]   _zz__30_14_inner_macOut_1;
  wire       [15:0]   _zz__30_14_inner_macOut_2;
  reg        [7:0]    _30_14_inner_activation;
  reg        [7:0]    _30_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_14_inner_macOut;

  assign _zz__zz__30_14_inner_macOut = ($signed(io_mulInput) * $signed(_30_14_inner_activation));
  assign _zz__zz__30_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_14_inner_macOut)) ? 16'h007f : _zz__30_14_inner_macOut_2);
  assign _zz__30_14_inner_macOut_2 = (($signed(_zz__30_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_14_inner_activation;
    end else begin
      io_macOut = _30_14_inner_macOut;
    end
  end

  assign _zz__30_14_inner_macOut = ($signed(_zz__zz__30_14_inner_macOut) + $signed(_zz__zz__30_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_14_inner_activation <= 8'h00;
      _30_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_14_inner_activation <= io_addInput;
      end else begin
        _30_14_inner_macOut <= _zz__30_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_973 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_13_inner_macOut;
  wire       [15:0]   _zz__zz__30_13_inner_macOut_1;
  wire       [15:0]   _zz__30_13_inner_macOut_1;
  wire       [15:0]   _zz__30_13_inner_macOut_2;
  reg        [7:0]    _30_13_inner_activation;
  reg        [7:0]    _30_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_13_inner_macOut;

  assign _zz__zz__30_13_inner_macOut = ($signed(io_mulInput) * $signed(_30_13_inner_activation));
  assign _zz__zz__30_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_13_inner_macOut)) ? 16'h007f : _zz__30_13_inner_macOut_2);
  assign _zz__30_13_inner_macOut_2 = (($signed(_zz__30_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_13_inner_activation;
    end else begin
      io_macOut = _30_13_inner_macOut;
    end
  end

  assign _zz__30_13_inner_macOut = ($signed(_zz__zz__30_13_inner_macOut) + $signed(_zz__zz__30_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_13_inner_activation <= 8'h00;
      _30_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_13_inner_activation <= io_addInput;
      end else begin
        _30_13_inner_macOut <= _zz__30_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_972 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_12_inner_macOut;
  wire       [15:0]   _zz__zz__30_12_inner_macOut_1;
  wire       [15:0]   _zz__30_12_inner_macOut_1;
  wire       [15:0]   _zz__30_12_inner_macOut_2;
  reg        [7:0]    _30_12_inner_activation;
  reg        [7:0]    _30_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_12_inner_macOut;

  assign _zz__zz__30_12_inner_macOut = ($signed(io_mulInput) * $signed(_30_12_inner_activation));
  assign _zz__zz__30_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_12_inner_macOut)) ? 16'h007f : _zz__30_12_inner_macOut_2);
  assign _zz__30_12_inner_macOut_2 = (($signed(_zz__30_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_12_inner_activation;
    end else begin
      io_macOut = _30_12_inner_macOut;
    end
  end

  assign _zz__30_12_inner_macOut = ($signed(_zz__zz__30_12_inner_macOut) + $signed(_zz__zz__30_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_12_inner_activation <= 8'h00;
      _30_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_12_inner_activation <= io_addInput;
      end else begin
        _30_12_inner_macOut <= _zz__30_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_971 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_11_inner_macOut;
  wire       [15:0]   _zz__zz__30_11_inner_macOut_1;
  wire       [15:0]   _zz__30_11_inner_macOut_1;
  wire       [15:0]   _zz__30_11_inner_macOut_2;
  reg        [7:0]    _30_11_inner_activation;
  reg        [7:0]    _30_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_11_inner_macOut;

  assign _zz__zz__30_11_inner_macOut = ($signed(io_mulInput) * $signed(_30_11_inner_activation));
  assign _zz__zz__30_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_11_inner_macOut)) ? 16'h007f : _zz__30_11_inner_macOut_2);
  assign _zz__30_11_inner_macOut_2 = (($signed(_zz__30_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_11_inner_activation;
    end else begin
      io_macOut = _30_11_inner_macOut;
    end
  end

  assign _zz__30_11_inner_macOut = ($signed(_zz__zz__30_11_inner_macOut) + $signed(_zz__zz__30_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_11_inner_activation <= 8'h00;
      _30_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_11_inner_activation <= io_addInput;
      end else begin
        _30_11_inner_macOut <= _zz__30_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_970 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_10_inner_macOut;
  wire       [15:0]   _zz__zz__30_10_inner_macOut_1;
  wire       [15:0]   _zz__30_10_inner_macOut_1;
  wire       [15:0]   _zz__30_10_inner_macOut_2;
  reg        [7:0]    _30_10_inner_activation;
  reg        [7:0]    _30_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_10_inner_macOut;

  assign _zz__zz__30_10_inner_macOut = ($signed(io_mulInput) * $signed(_30_10_inner_activation));
  assign _zz__zz__30_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_10_inner_macOut)) ? 16'h007f : _zz__30_10_inner_macOut_2);
  assign _zz__30_10_inner_macOut_2 = (($signed(_zz__30_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_10_inner_activation;
    end else begin
      io_macOut = _30_10_inner_macOut;
    end
  end

  assign _zz__30_10_inner_macOut = ($signed(_zz__zz__30_10_inner_macOut) + $signed(_zz__zz__30_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_10_inner_activation <= 8'h00;
      _30_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_10_inner_activation <= io_addInput;
      end else begin
        _30_10_inner_macOut <= _zz__30_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_969 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_9_inner_macOut;
  wire       [15:0]   _zz__zz__30_9_inner_macOut_1;
  wire       [15:0]   _zz__30_9_inner_macOut_1;
  wire       [15:0]   _zz__30_9_inner_macOut_2;
  reg        [7:0]    _30_9_inner_activation;
  reg        [7:0]    _30_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_9_inner_macOut;

  assign _zz__zz__30_9_inner_macOut = ($signed(io_mulInput) * $signed(_30_9_inner_activation));
  assign _zz__zz__30_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_9_inner_macOut)) ? 16'h007f : _zz__30_9_inner_macOut_2);
  assign _zz__30_9_inner_macOut_2 = (($signed(_zz__30_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_9_inner_activation;
    end else begin
      io_macOut = _30_9_inner_macOut;
    end
  end

  assign _zz__30_9_inner_macOut = ($signed(_zz__zz__30_9_inner_macOut) + $signed(_zz__zz__30_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_9_inner_activation <= 8'h00;
      _30_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_9_inner_activation <= io_addInput;
      end else begin
        _30_9_inner_macOut <= _zz__30_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_968 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_8_inner_macOut;
  wire       [15:0]   _zz__zz__30_8_inner_macOut_1;
  wire       [15:0]   _zz__30_8_inner_macOut_1;
  wire       [15:0]   _zz__30_8_inner_macOut_2;
  reg        [7:0]    _30_8_inner_activation;
  reg        [7:0]    _30_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_8_inner_macOut;

  assign _zz__zz__30_8_inner_macOut = ($signed(io_mulInput) * $signed(_30_8_inner_activation));
  assign _zz__zz__30_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_8_inner_macOut)) ? 16'h007f : _zz__30_8_inner_macOut_2);
  assign _zz__30_8_inner_macOut_2 = (($signed(_zz__30_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_8_inner_activation;
    end else begin
      io_macOut = _30_8_inner_macOut;
    end
  end

  assign _zz__30_8_inner_macOut = ($signed(_zz__zz__30_8_inner_macOut) + $signed(_zz__zz__30_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_8_inner_activation <= 8'h00;
      _30_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_8_inner_activation <= io_addInput;
      end else begin
        _30_8_inner_macOut <= _zz__30_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_967 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_7_inner_macOut;
  wire       [15:0]   _zz__zz__30_7_inner_macOut_1;
  wire       [15:0]   _zz__30_7_inner_macOut_1;
  wire       [15:0]   _zz__30_7_inner_macOut_2;
  reg        [7:0]    _30_7_inner_activation;
  reg        [7:0]    _30_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_7_inner_macOut;

  assign _zz__zz__30_7_inner_macOut = ($signed(io_mulInput) * $signed(_30_7_inner_activation));
  assign _zz__zz__30_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_7_inner_macOut)) ? 16'h007f : _zz__30_7_inner_macOut_2);
  assign _zz__30_7_inner_macOut_2 = (($signed(_zz__30_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_7_inner_activation;
    end else begin
      io_macOut = _30_7_inner_macOut;
    end
  end

  assign _zz__30_7_inner_macOut = ($signed(_zz__zz__30_7_inner_macOut) + $signed(_zz__zz__30_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_7_inner_activation <= 8'h00;
      _30_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_7_inner_activation <= io_addInput;
      end else begin
        _30_7_inner_macOut <= _zz__30_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_966 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_6_inner_macOut;
  wire       [15:0]   _zz__zz__30_6_inner_macOut_1;
  wire       [15:0]   _zz__30_6_inner_macOut_1;
  wire       [15:0]   _zz__30_6_inner_macOut_2;
  reg        [7:0]    _30_6_inner_activation;
  reg        [7:0]    _30_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_6_inner_macOut;

  assign _zz__zz__30_6_inner_macOut = ($signed(io_mulInput) * $signed(_30_6_inner_activation));
  assign _zz__zz__30_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_6_inner_macOut)) ? 16'h007f : _zz__30_6_inner_macOut_2);
  assign _zz__30_6_inner_macOut_2 = (($signed(_zz__30_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_6_inner_activation;
    end else begin
      io_macOut = _30_6_inner_macOut;
    end
  end

  assign _zz__30_6_inner_macOut = ($signed(_zz__zz__30_6_inner_macOut) + $signed(_zz__zz__30_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_6_inner_activation <= 8'h00;
      _30_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_6_inner_activation <= io_addInput;
      end else begin
        _30_6_inner_macOut <= _zz__30_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_965 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_5_inner_macOut;
  wire       [15:0]   _zz__zz__30_5_inner_macOut_1;
  wire       [15:0]   _zz__30_5_inner_macOut_1;
  wire       [15:0]   _zz__30_5_inner_macOut_2;
  reg        [7:0]    _30_5_inner_activation;
  reg        [7:0]    _30_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_5_inner_macOut;

  assign _zz__zz__30_5_inner_macOut = ($signed(io_mulInput) * $signed(_30_5_inner_activation));
  assign _zz__zz__30_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_5_inner_macOut)) ? 16'h007f : _zz__30_5_inner_macOut_2);
  assign _zz__30_5_inner_macOut_2 = (($signed(_zz__30_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_5_inner_activation;
    end else begin
      io_macOut = _30_5_inner_macOut;
    end
  end

  assign _zz__30_5_inner_macOut = ($signed(_zz__zz__30_5_inner_macOut) + $signed(_zz__zz__30_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_5_inner_activation <= 8'h00;
      _30_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_5_inner_activation <= io_addInput;
      end else begin
        _30_5_inner_macOut <= _zz__30_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_964 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_4_inner_macOut;
  wire       [15:0]   _zz__zz__30_4_inner_macOut_1;
  wire       [15:0]   _zz__30_4_inner_macOut_1;
  wire       [15:0]   _zz__30_4_inner_macOut_2;
  reg        [7:0]    _30_4_inner_activation;
  reg        [7:0]    _30_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_4_inner_macOut;

  assign _zz__zz__30_4_inner_macOut = ($signed(io_mulInput) * $signed(_30_4_inner_activation));
  assign _zz__zz__30_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_4_inner_macOut)) ? 16'h007f : _zz__30_4_inner_macOut_2);
  assign _zz__30_4_inner_macOut_2 = (($signed(_zz__30_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_4_inner_activation;
    end else begin
      io_macOut = _30_4_inner_macOut;
    end
  end

  assign _zz__30_4_inner_macOut = ($signed(_zz__zz__30_4_inner_macOut) + $signed(_zz__zz__30_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_4_inner_activation <= 8'h00;
      _30_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_4_inner_activation <= io_addInput;
      end else begin
        _30_4_inner_macOut <= _zz__30_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_963 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_3_inner_macOut;
  wire       [15:0]   _zz__zz__30_3_inner_macOut_1;
  wire       [15:0]   _zz__30_3_inner_macOut_1;
  wire       [15:0]   _zz__30_3_inner_macOut_2;
  reg        [7:0]    _30_3_inner_activation;
  reg        [7:0]    _30_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_3_inner_macOut;

  assign _zz__zz__30_3_inner_macOut = ($signed(io_mulInput) * $signed(_30_3_inner_activation));
  assign _zz__zz__30_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_3_inner_macOut)) ? 16'h007f : _zz__30_3_inner_macOut_2);
  assign _zz__30_3_inner_macOut_2 = (($signed(_zz__30_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_3_inner_activation;
    end else begin
      io_macOut = _30_3_inner_macOut;
    end
  end

  assign _zz__30_3_inner_macOut = ($signed(_zz__zz__30_3_inner_macOut) + $signed(_zz__zz__30_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_3_inner_activation <= 8'h00;
      _30_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_3_inner_activation <= io_addInput;
      end else begin
        _30_3_inner_macOut <= _zz__30_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_962 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_2_inner_macOut;
  wire       [15:0]   _zz__zz__30_2_inner_macOut_1;
  wire       [15:0]   _zz__30_2_inner_macOut_1;
  wire       [15:0]   _zz__30_2_inner_macOut_2;
  reg        [7:0]    _30_2_inner_activation;
  reg        [7:0]    _30_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_2_inner_macOut;

  assign _zz__zz__30_2_inner_macOut = ($signed(io_mulInput) * $signed(_30_2_inner_activation));
  assign _zz__zz__30_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_2_inner_macOut)) ? 16'h007f : _zz__30_2_inner_macOut_2);
  assign _zz__30_2_inner_macOut_2 = (($signed(_zz__30_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_2_inner_activation;
    end else begin
      io_macOut = _30_2_inner_macOut;
    end
  end

  assign _zz__30_2_inner_macOut = ($signed(_zz__zz__30_2_inner_macOut) + $signed(_zz__zz__30_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_2_inner_activation <= 8'h00;
      _30_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_2_inner_activation <= io_addInput;
      end else begin
        _30_2_inner_macOut <= _zz__30_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_961 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_1_inner_macOut;
  wire       [15:0]   _zz__zz__30_1_inner_macOut_1;
  wire       [15:0]   _zz__30_1_inner_macOut_1;
  wire       [15:0]   _zz__30_1_inner_macOut_2;
  reg        [7:0]    _30_1_inner_activation;
  reg        [7:0]    _30_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_1_inner_macOut;

  assign _zz__zz__30_1_inner_macOut = ($signed(io_mulInput) * $signed(_30_1_inner_activation));
  assign _zz__zz__30_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_1_inner_macOut)) ? 16'h007f : _zz__30_1_inner_macOut_2);
  assign _zz__30_1_inner_macOut_2 = (($signed(_zz__30_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_1_inner_activation;
    end else begin
      io_macOut = _30_1_inner_macOut;
    end
  end

  assign _zz__30_1_inner_macOut = ($signed(_zz__zz__30_1_inner_macOut) + $signed(_zz__zz__30_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_1_inner_activation <= 8'h00;
      _30_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_1_inner_activation <= io_addInput;
      end else begin
        _30_1_inner_macOut <= _zz__30_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_960 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__30_0_inner_macOut;
  wire       [15:0]   _zz__zz__30_0_inner_macOut_1;
  wire       [15:0]   _zz__30_0_inner_macOut_1;
  wire       [15:0]   _zz__30_0_inner_macOut_2;
  reg        [7:0]    _30_0_inner_activation;
  reg        [7:0]    _30_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__30_0_inner_macOut;

  assign _zz__zz__30_0_inner_macOut = ($signed(io_mulInput) * $signed(_30_0_inner_activation));
  assign _zz__zz__30_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__30_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__30_0_inner_macOut)) ? 16'h007f : _zz__30_0_inner_macOut_2);
  assign _zz__30_0_inner_macOut_2 = (($signed(_zz__30_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__30_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _30_0_inner_activation;
    end else begin
      io_macOut = _30_0_inner_macOut;
    end
  end

  assign _zz__30_0_inner_macOut = ($signed(_zz__zz__30_0_inner_macOut) + $signed(_zz__zz__30_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _30_0_inner_activation <= 8'h00;
      _30_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _30_0_inner_activation <= io_addInput;
      end else begin
        _30_0_inner_macOut <= _zz__30_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_959 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_31_inner_macOut;
  wire       [15:0]   _zz__zz__29_31_inner_macOut_1;
  wire       [15:0]   _zz__29_31_inner_macOut_1;
  wire       [15:0]   _zz__29_31_inner_macOut_2;
  reg        [7:0]    _29_31_inner_activation;
  reg        [7:0]    _29_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_31_inner_macOut;

  assign _zz__zz__29_31_inner_macOut = ($signed(io_mulInput) * $signed(_29_31_inner_activation));
  assign _zz__zz__29_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_31_inner_macOut)) ? 16'h007f : _zz__29_31_inner_macOut_2);
  assign _zz__29_31_inner_macOut_2 = (($signed(_zz__29_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_31_inner_activation;
    end else begin
      io_macOut = _29_31_inner_macOut;
    end
  end

  assign _zz__29_31_inner_macOut = ($signed(_zz__zz__29_31_inner_macOut) + $signed(_zz__zz__29_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_31_inner_activation <= 8'h00;
      _29_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_31_inner_activation <= io_addInput;
      end else begin
        _29_31_inner_macOut <= _zz__29_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_958 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_30_inner_macOut;
  wire       [15:0]   _zz__zz__29_30_inner_macOut_1;
  wire       [15:0]   _zz__29_30_inner_macOut_1;
  wire       [15:0]   _zz__29_30_inner_macOut_2;
  reg        [7:0]    _29_30_inner_activation;
  reg        [7:0]    _29_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_30_inner_macOut;

  assign _zz__zz__29_30_inner_macOut = ($signed(io_mulInput) * $signed(_29_30_inner_activation));
  assign _zz__zz__29_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_30_inner_macOut)) ? 16'h007f : _zz__29_30_inner_macOut_2);
  assign _zz__29_30_inner_macOut_2 = (($signed(_zz__29_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_30_inner_activation;
    end else begin
      io_macOut = _29_30_inner_macOut;
    end
  end

  assign _zz__29_30_inner_macOut = ($signed(_zz__zz__29_30_inner_macOut) + $signed(_zz__zz__29_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_30_inner_activation <= 8'h00;
      _29_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_30_inner_activation <= io_addInput;
      end else begin
        _29_30_inner_macOut <= _zz__29_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_957 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_29_inner_macOut;
  wire       [15:0]   _zz__zz__29_29_inner_macOut_1;
  wire       [15:0]   _zz__29_29_inner_macOut_1;
  wire       [15:0]   _zz__29_29_inner_macOut_2;
  reg        [7:0]    _29_29_inner_activation;
  reg        [7:0]    _29_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_29_inner_macOut;

  assign _zz__zz__29_29_inner_macOut = ($signed(io_mulInput) * $signed(_29_29_inner_activation));
  assign _zz__zz__29_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_29_inner_macOut)) ? 16'h007f : _zz__29_29_inner_macOut_2);
  assign _zz__29_29_inner_macOut_2 = (($signed(_zz__29_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_29_inner_activation;
    end else begin
      io_macOut = _29_29_inner_macOut;
    end
  end

  assign _zz__29_29_inner_macOut = ($signed(_zz__zz__29_29_inner_macOut) + $signed(_zz__zz__29_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_29_inner_activation <= 8'h00;
      _29_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_29_inner_activation <= io_addInput;
      end else begin
        _29_29_inner_macOut <= _zz__29_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_956 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_28_inner_macOut;
  wire       [15:0]   _zz__zz__29_28_inner_macOut_1;
  wire       [15:0]   _zz__29_28_inner_macOut_1;
  wire       [15:0]   _zz__29_28_inner_macOut_2;
  reg        [7:0]    _29_28_inner_activation;
  reg        [7:0]    _29_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_28_inner_macOut;

  assign _zz__zz__29_28_inner_macOut = ($signed(io_mulInput) * $signed(_29_28_inner_activation));
  assign _zz__zz__29_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_28_inner_macOut)) ? 16'h007f : _zz__29_28_inner_macOut_2);
  assign _zz__29_28_inner_macOut_2 = (($signed(_zz__29_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_28_inner_activation;
    end else begin
      io_macOut = _29_28_inner_macOut;
    end
  end

  assign _zz__29_28_inner_macOut = ($signed(_zz__zz__29_28_inner_macOut) + $signed(_zz__zz__29_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_28_inner_activation <= 8'h00;
      _29_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_28_inner_activation <= io_addInput;
      end else begin
        _29_28_inner_macOut <= _zz__29_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_955 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_27_inner_macOut;
  wire       [15:0]   _zz__zz__29_27_inner_macOut_1;
  wire       [15:0]   _zz__29_27_inner_macOut_1;
  wire       [15:0]   _zz__29_27_inner_macOut_2;
  reg        [7:0]    _29_27_inner_activation;
  reg        [7:0]    _29_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_27_inner_macOut;

  assign _zz__zz__29_27_inner_macOut = ($signed(io_mulInput) * $signed(_29_27_inner_activation));
  assign _zz__zz__29_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_27_inner_macOut)) ? 16'h007f : _zz__29_27_inner_macOut_2);
  assign _zz__29_27_inner_macOut_2 = (($signed(_zz__29_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_27_inner_activation;
    end else begin
      io_macOut = _29_27_inner_macOut;
    end
  end

  assign _zz__29_27_inner_macOut = ($signed(_zz__zz__29_27_inner_macOut) + $signed(_zz__zz__29_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_27_inner_activation <= 8'h00;
      _29_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_27_inner_activation <= io_addInput;
      end else begin
        _29_27_inner_macOut <= _zz__29_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_954 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_26_inner_macOut;
  wire       [15:0]   _zz__zz__29_26_inner_macOut_1;
  wire       [15:0]   _zz__29_26_inner_macOut_1;
  wire       [15:0]   _zz__29_26_inner_macOut_2;
  reg        [7:0]    _29_26_inner_activation;
  reg        [7:0]    _29_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_26_inner_macOut;

  assign _zz__zz__29_26_inner_macOut = ($signed(io_mulInput) * $signed(_29_26_inner_activation));
  assign _zz__zz__29_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_26_inner_macOut)) ? 16'h007f : _zz__29_26_inner_macOut_2);
  assign _zz__29_26_inner_macOut_2 = (($signed(_zz__29_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_26_inner_activation;
    end else begin
      io_macOut = _29_26_inner_macOut;
    end
  end

  assign _zz__29_26_inner_macOut = ($signed(_zz__zz__29_26_inner_macOut) + $signed(_zz__zz__29_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_26_inner_activation <= 8'h00;
      _29_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_26_inner_activation <= io_addInput;
      end else begin
        _29_26_inner_macOut <= _zz__29_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_953 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_25_inner_macOut;
  wire       [15:0]   _zz__zz__29_25_inner_macOut_1;
  wire       [15:0]   _zz__29_25_inner_macOut_1;
  wire       [15:0]   _zz__29_25_inner_macOut_2;
  reg        [7:0]    _29_25_inner_activation;
  reg        [7:0]    _29_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_25_inner_macOut;

  assign _zz__zz__29_25_inner_macOut = ($signed(io_mulInput) * $signed(_29_25_inner_activation));
  assign _zz__zz__29_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_25_inner_macOut)) ? 16'h007f : _zz__29_25_inner_macOut_2);
  assign _zz__29_25_inner_macOut_2 = (($signed(_zz__29_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_25_inner_activation;
    end else begin
      io_macOut = _29_25_inner_macOut;
    end
  end

  assign _zz__29_25_inner_macOut = ($signed(_zz__zz__29_25_inner_macOut) + $signed(_zz__zz__29_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_25_inner_activation <= 8'h00;
      _29_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_25_inner_activation <= io_addInput;
      end else begin
        _29_25_inner_macOut <= _zz__29_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_952 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_24_inner_macOut;
  wire       [15:0]   _zz__zz__29_24_inner_macOut_1;
  wire       [15:0]   _zz__29_24_inner_macOut_1;
  wire       [15:0]   _zz__29_24_inner_macOut_2;
  reg        [7:0]    _29_24_inner_activation;
  reg        [7:0]    _29_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_24_inner_macOut;

  assign _zz__zz__29_24_inner_macOut = ($signed(io_mulInput) * $signed(_29_24_inner_activation));
  assign _zz__zz__29_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_24_inner_macOut)) ? 16'h007f : _zz__29_24_inner_macOut_2);
  assign _zz__29_24_inner_macOut_2 = (($signed(_zz__29_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_24_inner_activation;
    end else begin
      io_macOut = _29_24_inner_macOut;
    end
  end

  assign _zz__29_24_inner_macOut = ($signed(_zz__zz__29_24_inner_macOut) + $signed(_zz__zz__29_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_24_inner_activation <= 8'h00;
      _29_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_24_inner_activation <= io_addInput;
      end else begin
        _29_24_inner_macOut <= _zz__29_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_951 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_23_inner_macOut;
  wire       [15:0]   _zz__zz__29_23_inner_macOut_1;
  wire       [15:0]   _zz__29_23_inner_macOut_1;
  wire       [15:0]   _zz__29_23_inner_macOut_2;
  reg        [7:0]    _29_23_inner_activation;
  reg        [7:0]    _29_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_23_inner_macOut;

  assign _zz__zz__29_23_inner_macOut = ($signed(io_mulInput) * $signed(_29_23_inner_activation));
  assign _zz__zz__29_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_23_inner_macOut)) ? 16'h007f : _zz__29_23_inner_macOut_2);
  assign _zz__29_23_inner_macOut_2 = (($signed(_zz__29_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_23_inner_activation;
    end else begin
      io_macOut = _29_23_inner_macOut;
    end
  end

  assign _zz__29_23_inner_macOut = ($signed(_zz__zz__29_23_inner_macOut) + $signed(_zz__zz__29_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_23_inner_activation <= 8'h00;
      _29_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_23_inner_activation <= io_addInput;
      end else begin
        _29_23_inner_macOut <= _zz__29_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_950 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_22_inner_macOut;
  wire       [15:0]   _zz__zz__29_22_inner_macOut_1;
  wire       [15:0]   _zz__29_22_inner_macOut_1;
  wire       [15:0]   _zz__29_22_inner_macOut_2;
  reg        [7:0]    _29_22_inner_activation;
  reg        [7:0]    _29_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_22_inner_macOut;

  assign _zz__zz__29_22_inner_macOut = ($signed(io_mulInput) * $signed(_29_22_inner_activation));
  assign _zz__zz__29_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_22_inner_macOut)) ? 16'h007f : _zz__29_22_inner_macOut_2);
  assign _zz__29_22_inner_macOut_2 = (($signed(_zz__29_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_22_inner_activation;
    end else begin
      io_macOut = _29_22_inner_macOut;
    end
  end

  assign _zz__29_22_inner_macOut = ($signed(_zz__zz__29_22_inner_macOut) + $signed(_zz__zz__29_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_22_inner_activation <= 8'h00;
      _29_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_22_inner_activation <= io_addInput;
      end else begin
        _29_22_inner_macOut <= _zz__29_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_949 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_21_inner_macOut;
  wire       [15:0]   _zz__zz__29_21_inner_macOut_1;
  wire       [15:0]   _zz__29_21_inner_macOut_1;
  wire       [15:0]   _zz__29_21_inner_macOut_2;
  reg        [7:0]    _29_21_inner_activation;
  reg        [7:0]    _29_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_21_inner_macOut;

  assign _zz__zz__29_21_inner_macOut = ($signed(io_mulInput) * $signed(_29_21_inner_activation));
  assign _zz__zz__29_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_21_inner_macOut)) ? 16'h007f : _zz__29_21_inner_macOut_2);
  assign _zz__29_21_inner_macOut_2 = (($signed(_zz__29_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_21_inner_activation;
    end else begin
      io_macOut = _29_21_inner_macOut;
    end
  end

  assign _zz__29_21_inner_macOut = ($signed(_zz__zz__29_21_inner_macOut) + $signed(_zz__zz__29_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_21_inner_activation <= 8'h00;
      _29_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_21_inner_activation <= io_addInput;
      end else begin
        _29_21_inner_macOut <= _zz__29_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_948 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_20_inner_macOut;
  wire       [15:0]   _zz__zz__29_20_inner_macOut_1;
  wire       [15:0]   _zz__29_20_inner_macOut_1;
  wire       [15:0]   _zz__29_20_inner_macOut_2;
  reg        [7:0]    _29_20_inner_activation;
  reg        [7:0]    _29_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_20_inner_macOut;

  assign _zz__zz__29_20_inner_macOut = ($signed(io_mulInput) * $signed(_29_20_inner_activation));
  assign _zz__zz__29_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_20_inner_macOut)) ? 16'h007f : _zz__29_20_inner_macOut_2);
  assign _zz__29_20_inner_macOut_2 = (($signed(_zz__29_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_20_inner_activation;
    end else begin
      io_macOut = _29_20_inner_macOut;
    end
  end

  assign _zz__29_20_inner_macOut = ($signed(_zz__zz__29_20_inner_macOut) + $signed(_zz__zz__29_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_20_inner_activation <= 8'h00;
      _29_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_20_inner_activation <= io_addInput;
      end else begin
        _29_20_inner_macOut <= _zz__29_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_947 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_19_inner_macOut;
  wire       [15:0]   _zz__zz__29_19_inner_macOut_1;
  wire       [15:0]   _zz__29_19_inner_macOut_1;
  wire       [15:0]   _zz__29_19_inner_macOut_2;
  reg        [7:0]    _29_19_inner_activation;
  reg        [7:0]    _29_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_19_inner_macOut;

  assign _zz__zz__29_19_inner_macOut = ($signed(io_mulInput) * $signed(_29_19_inner_activation));
  assign _zz__zz__29_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_19_inner_macOut)) ? 16'h007f : _zz__29_19_inner_macOut_2);
  assign _zz__29_19_inner_macOut_2 = (($signed(_zz__29_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_19_inner_activation;
    end else begin
      io_macOut = _29_19_inner_macOut;
    end
  end

  assign _zz__29_19_inner_macOut = ($signed(_zz__zz__29_19_inner_macOut) + $signed(_zz__zz__29_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_19_inner_activation <= 8'h00;
      _29_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_19_inner_activation <= io_addInput;
      end else begin
        _29_19_inner_macOut <= _zz__29_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_946 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_18_inner_macOut;
  wire       [15:0]   _zz__zz__29_18_inner_macOut_1;
  wire       [15:0]   _zz__29_18_inner_macOut_1;
  wire       [15:0]   _zz__29_18_inner_macOut_2;
  reg        [7:0]    _29_18_inner_activation;
  reg        [7:0]    _29_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_18_inner_macOut;

  assign _zz__zz__29_18_inner_macOut = ($signed(io_mulInput) * $signed(_29_18_inner_activation));
  assign _zz__zz__29_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_18_inner_macOut)) ? 16'h007f : _zz__29_18_inner_macOut_2);
  assign _zz__29_18_inner_macOut_2 = (($signed(_zz__29_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_18_inner_activation;
    end else begin
      io_macOut = _29_18_inner_macOut;
    end
  end

  assign _zz__29_18_inner_macOut = ($signed(_zz__zz__29_18_inner_macOut) + $signed(_zz__zz__29_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_18_inner_activation <= 8'h00;
      _29_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_18_inner_activation <= io_addInput;
      end else begin
        _29_18_inner_macOut <= _zz__29_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_945 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_17_inner_macOut;
  wire       [15:0]   _zz__zz__29_17_inner_macOut_1;
  wire       [15:0]   _zz__29_17_inner_macOut_1;
  wire       [15:0]   _zz__29_17_inner_macOut_2;
  reg        [7:0]    _29_17_inner_activation;
  reg        [7:0]    _29_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_17_inner_macOut;

  assign _zz__zz__29_17_inner_macOut = ($signed(io_mulInput) * $signed(_29_17_inner_activation));
  assign _zz__zz__29_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_17_inner_macOut)) ? 16'h007f : _zz__29_17_inner_macOut_2);
  assign _zz__29_17_inner_macOut_2 = (($signed(_zz__29_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_17_inner_activation;
    end else begin
      io_macOut = _29_17_inner_macOut;
    end
  end

  assign _zz__29_17_inner_macOut = ($signed(_zz__zz__29_17_inner_macOut) + $signed(_zz__zz__29_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_17_inner_activation <= 8'h00;
      _29_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_17_inner_activation <= io_addInput;
      end else begin
        _29_17_inner_macOut <= _zz__29_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_944 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_16_inner_macOut;
  wire       [15:0]   _zz__zz__29_16_inner_macOut_1;
  wire       [15:0]   _zz__29_16_inner_macOut_1;
  wire       [15:0]   _zz__29_16_inner_macOut_2;
  reg        [7:0]    _29_16_inner_activation;
  reg        [7:0]    _29_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_16_inner_macOut;

  assign _zz__zz__29_16_inner_macOut = ($signed(io_mulInput) * $signed(_29_16_inner_activation));
  assign _zz__zz__29_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_16_inner_macOut)) ? 16'h007f : _zz__29_16_inner_macOut_2);
  assign _zz__29_16_inner_macOut_2 = (($signed(_zz__29_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_16_inner_activation;
    end else begin
      io_macOut = _29_16_inner_macOut;
    end
  end

  assign _zz__29_16_inner_macOut = ($signed(_zz__zz__29_16_inner_macOut) + $signed(_zz__zz__29_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_16_inner_activation <= 8'h00;
      _29_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_16_inner_activation <= io_addInput;
      end else begin
        _29_16_inner_macOut <= _zz__29_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_943 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_15_inner_macOut;
  wire       [15:0]   _zz__zz__29_15_inner_macOut_1;
  wire       [15:0]   _zz__29_15_inner_macOut_1;
  wire       [15:0]   _zz__29_15_inner_macOut_2;
  reg        [7:0]    _29_15_inner_activation;
  reg        [7:0]    _29_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_15_inner_macOut;

  assign _zz__zz__29_15_inner_macOut = ($signed(io_mulInput) * $signed(_29_15_inner_activation));
  assign _zz__zz__29_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_15_inner_macOut)) ? 16'h007f : _zz__29_15_inner_macOut_2);
  assign _zz__29_15_inner_macOut_2 = (($signed(_zz__29_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_15_inner_activation;
    end else begin
      io_macOut = _29_15_inner_macOut;
    end
  end

  assign _zz__29_15_inner_macOut = ($signed(_zz__zz__29_15_inner_macOut) + $signed(_zz__zz__29_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_15_inner_activation <= 8'h00;
      _29_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_15_inner_activation <= io_addInput;
      end else begin
        _29_15_inner_macOut <= _zz__29_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_942 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_14_inner_macOut;
  wire       [15:0]   _zz__zz__29_14_inner_macOut_1;
  wire       [15:0]   _zz__29_14_inner_macOut_1;
  wire       [15:0]   _zz__29_14_inner_macOut_2;
  reg        [7:0]    _29_14_inner_activation;
  reg        [7:0]    _29_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_14_inner_macOut;

  assign _zz__zz__29_14_inner_macOut = ($signed(io_mulInput) * $signed(_29_14_inner_activation));
  assign _zz__zz__29_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_14_inner_macOut)) ? 16'h007f : _zz__29_14_inner_macOut_2);
  assign _zz__29_14_inner_macOut_2 = (($signed(_zz__29_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_14_inner_activation;
    end else begin
      io_macOut = _29_14_inner_macOut;
    end
  end

  assign _zz__29_14_inner_macOut = ($signed(_zz__zz__29_14_inner_macOut) + $signed(_zz__zz__29_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_14_inner_activation <= 8'h00;
      _29_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_14_inner_activation <= io_addInput;
      end else begin
        _29_14_inner_macOut <= _zz__29_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_941 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_13_inner_macOut;
  wire       [15:0]   _zz__zz__29_13_inner_macOut_1;
  wire       [15:0]   _zz__29_13_inner_macOut_1;
  wire       [15:0]   _zz__29_13_inner_macOut_2;
  reg        [7:0]    _29_13_inner_activation;
  reg        [7:0]    _29_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_13_inner_macOut;

  assign _zz__zz__29_13_inner_macOut = ($signed(io_mulInput) * $signed(_29_13_inner_activation));
  assign _zz__zz__29_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_13_inner_macOut)) ? 16'h007f : _zz__29_13_inner_macOut_2);
  assign _zz__29_13_inner_macOut_2 = (($signed(_zz__29_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_13_inner_activation;
    end else begin
      io_macOut = _29_13_inner_macOut;
    end
  end

  assign _zz__29_13_inner_macOut = ($signed(_zz__zz__29_13_inner_macOut) + $signed(_zz__zz__29_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_13_inner_activation <= 8'h00;
      _29_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_13_inner_activation <= io_addInput;
      end else begin
        _29_13_inner_macOut <= _zz__29_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_940 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_12_inner_macOut;
  wire       [15:0]   _zz__zz__29_12_inner_macOut_1;
  wire       [15:0]   _zz__29_12_inner_macOut_1;
  wire       [15:0]   _zz__29_12_inner_macOut_2;
  reg        [7:0]    _29_12_inner_activation;
  reg        [7:0]    _29_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_12_inner_macOut;

  assign _zz__zz__29_12_inner_macOut = ($signed(io_mulInput) * $signed(_29_12_inner_activation));
  assign _zz__zz__29_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_12_inner_macOut)) ? 16'h007f : _zz__29_12_inner_macOut_2);
  assign _zz__29_12_inner_macOut_2 = (($signed(_zz__29_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_12_inner_activation;
    end else begin
      io_macOut = _29_12_inner_macOut;
    end
  end

  assign _zz__29_12_inner_macOut = ($signed(_zz__zz__29_12_inner_macOut) + $signed(_zz__zz__29_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_12_inner_activation <= 8'h00;
      _29_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_12_inner_activation <= io_addInput;
      end else begin
        _29_12_inner_macOut <= _zz__29_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_939 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_11_inner_macOut;
  wire       [15:0]   _zz__zz__29_11_inner_macOut_1;
  wire       [15:0]   _zz__29_11_inner_macOut_1;
  wire       [15:0]   _zz__29_11_inner_macOut_2;
  reg        [7:0]    _29_11_inner_activation;
  reg        [7:0]    _29_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_11_inner_macOut;

  assign _zz__zz__29_11_inner_macOut = ($signed(io_mulInput) * $signed(_29_11_inner_activation));
  assign _zz__zz__29_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_11_inner_macOut)) ? 16'h007f : _zz__29_11_inner_macOut_2);
  assign _zz__29_11_inner_macOut_2 = (($signed(_zz__29_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_11_inner_activation;
    end else begin
      io_macOut = _29_11_inner_macOut;
    end
  end

  assign _zz__29_11_inner_macOut = ($signed(_zz__zz__29_11_inner_macOut) + $signed(_zz__zz__29_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_11_inner_activation <= 8'h00;
      _29_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_11_inner_activation <= io_addInput;
      end else begin
        _29_11_inner_macOut <= _zz__29_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_938 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_10_inner_macOut;
  wire       [15:0]   _zz__zz__29_10_inner_macOut_1;
  wire       [15:0]   _zz__29_10_inner_macOut_1;
  wire       [15:0]   _zz__29_10_inner_macOut_2;
  reg        [7:0]    _29_10_inner_activation;
  reg        [7:0]    _29_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_10_inner_macOut;

  assign _zz__zz__29_10_inner_macOut = ($signed(io_mulInput) * $signed(_29_10_inner_activation));
  assign _zz__zz__29_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_10_inner_macOut)) ? 16'h007f : _zz__29_10_inner_macOut_2);
  assign _zz__29_10_inner_macOut_2 = (($signed(_zz__29_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_10_inner_activation;
    end else begin
      io_macOut = _29_10_inner_macOut;
    end
  end

  assign _zz__29_10_inner_macOut = ($signed(_zz__zz__29_10_inner_macOut) + $signed(_zz__zz__29_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_10_inner_activation <= 8'h00;
      _29_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_10_inner_activation <= io_addInput;
      end else begin
        _29_10_inner_macOut <= _zz__29_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_937 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_9_inner_macOut;
  wire       [15:0]   _zz__zz__29_9_inner_macOut_1;
  wire       [15:0]   _zz__29_9_inner_macOut_1;
  wire       [15:0]   _zz__29_9_inner_macOut_2;
  reg        [7:0]    _29_9_inner_activation;
  reg        [7:0]    _29_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_9_inner_macOut;

  assign _zz__zz__29_9_inner_macOut = ($signed(io_mulInput) * $signed(_29_9_inner_activation));
  assign _zz__zz__29_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_9_inner_macOut)) ? 16'h007f : _zz__29_9_inner_macOut_2);
  assign _zz__29_9_inner_macOut_2 = (($signed(_zz__29_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_9_inner_activation;
    end else begin
      io_macOut = _29_9_inner_macOut;
    end
  end

  assign _zz__29_9_inner_macOut = ($signed(_zz__zz__29_9_inner_macOut) + $signed(_zz__zz__29_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_9_inner_activation <= 8'h00;
      _29_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_9_inner_activation <= io_addInput;
      end else begin
        _29_9_inner_macOut <= _zz__29_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_936 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_8_inner_macOut;
  wire       [15:0]   _zz__zz__29_8_inner_macOut_1;
  wire       [15:0]   _zz__29_8_inner_macOut_1;
  wire       [15:0]   _zz__29_8_inner_macOut_2;
  reg        [7:0]    _29_8_inner_activation;
  reg        [7:0]    _29_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_8_inner_macOut;

  assign _zz__zz__29_8_inner_macOut = ($signed(io_mulInput) * $signed(_29_8_inner_activation));
  assign _zz__zz__29_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_8_inner_macOut)) ? 16'h007f : _zz__29_8_inner_macOut_2);
  assign _zz__29_8_inner_macOut_2 = (($signed(_zz__29_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_8_inner_activation;
    end else begin
      io_macOut = _29_8_inner_macOut;
    end
  end

  assign _zz__29_8_inner_macOut = ($signed(_zz__zz__29_8_inner_macOut) + $signed(_zz__zz__29_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_8_inner_activation <= 8'h00;
      _29_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_8_inner_activation <= io_addInput;
      end else begin
        _29_8_inner_macOut <= _zz__29_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_935 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_7_inner_macOut;
  wire       [15:0]   _zz__zz__29_7_inner_macOut_1;
  wire       [15:0]   _zz__29_7_inner_macOut_1;
  wire       [15:0]   _zz__29_7_inner_macOut_2;
  reg        [7:0]    _29_7_inner_activation;
  reg        [7:0]    _29_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_7_inner_macOut;

  assign _zz__zz__29_7_inner_macOut = ($signed(io_mulInput) * $signed(_29_7_inner_activation));
  assign _zz__zz__29_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_7_inner_macOut)) ? 16'h007f : _zz__29_7_inner_macOut_2);
  assign _zz__29_7_inner_macOut_2 = (($signed(_zz__29_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_7_inner_activation;
    end else begin
      io_macOut = _29_7_inner_macOut;
    end
  end

  assign _zz__29_7_inner_macOut = ($signed(_zz__zz__29_7_inner_macOut) + $signed(_zz__zz__29_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_7_inner_activation <= 8'h00;
      _29_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_7_inner_activation <= io_addInput;
      end else begin
        _29_7_inner_macOut <= _zz__29_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_934 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_6_inner_macOut;
  wire       [15:0]   _zz__zz__29_6_inner_macOut_1;
  wire       [15:0]   _zz__29_6_inner_macOut_1;
  wire       [15:0]   _zz__29_6_inner_macOut_2;
  reg        [7:0]    _29_6_inner_activation;
  reg        [7:0]    _29_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_6_inner_macOut;

  assign _zz__zz__29_6_inner_macOut = ($signed(io_mulInput) * $signed(_29_6_inner_activation));
  assign _zz__zz__29_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_6_inner_macOut)) ? 16'h007f : _zz__29_6_inner_macOut_2);
  assign _zz__29_6_inner_macOut_2 = (($signed(_zz__29_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_6_inner_activation;
    end else begin
      io_macOut = _29_6_inner_macOut;
    end
  end

  assign _zz__29_6_inner_macOut = ($signed(_zz__zz__29_6_inner_macOut) + $signed(_zz__zz__29_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_6_inner_activation <= 8'h00;
      _29_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_6_inner_activation <= io_addInput;
      end else begin
        _29_6_inner_macOut <= _zz__29_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_933 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_5_inner_macOut;
  wire       [15:0]   _zz__zz__29_5_inner_macOut_1;
  wire       [15:0]   _zz__29_5_inner_macOut_1;
  wire       [15:0]   _zz__29_5_inner_macOut_2;
  reg        [7:0]    _29_5_inner_activation;
  reg        [7:0]    _29_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_5_inner_macOut;

  assign _zz__zz__29_5_inner_macOut = ($signed(io_mulInput) * $signed(_29_5_inner_activation));
  assign _zz__zz__29_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_5_inner_macOut)) ? 16'h007f : _zz__29_5_inner_macOut_2);
  assign _zz__29_5_inner_macOut_2 = (($signed(_zz__29_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_5_inner_activation;
    end else begin
      io_macOut = _29_5_inner_macOut;
    end
  end

  assign _zz__29_5_inner_macOut = ($signed(_zz__zz__29_5_inner_macOut) + $signed(_zz__zz__29_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_5_inner_activation <= 8'h00;
      _29_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_5_inner_activation <= io_addInput;
      end else begin
        _29_5_inner_macOut <= _zz__29_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_932 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_4_inner_macOut;
  wire       [15:0]   _zz__zz__29_4_inner_macOut_1;
  wire       [15:0]   _zz__29_4_inner_macOut_1;
  wire       [15:0]   _zz__29_4_inner_macOut_2;
  reg        [7:0]    _29_4_inner_activation;
  reg        [7:0]    _29_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_4_inner_macOut;

  assign _zz__zz__29_4_inner_macOut = ($signed(io_mulInput) * $signed(_29_4_inner_activation));
  assign _zz__zz__29_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_4_inner_macOut)) ? 16'h007f : _zz__29_4_inner_macOut_2);
  assign _zz__29_4_inner_macOut_2 = (($signed(_zz__29_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_4_inner_activation;
    end else begin
      io_macOut = _29_4_inner_macOut;
    end
  end

  assign _zz__29_4_inner_macOut = ($signed(_zz__zz__29_4_inner_macOut) + $signed(_zz__zz__29_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_4_inner_activation <= 8'h00;
      _29_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_4_inner_activation <= io_addInput;
      end else begin
        _29_4_inner_macOut <= _zz__29_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_931 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_3_inner_macOut;
  wire       [15:0]   _zz__zz__29_3_inner_macOut_1;
  wire       [15:0]   _zz__29_3_inner_macOut_1;
  wire       [15:0]   _zz__29_3_inner_macOut_2;
  reg        [7:0]    _29_3_inner_activation;
  reg        [7:0]    _29_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_3_inner_macOut;

  assign _zz__zz__29_3_inner_macOut = ($signed(io_mulInput) * $signed(_29_3_inner_activation));
  assign _zz__zz__29_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_3_inner_macOut)) ? 16'h007f : _zz__29_3_inner_macOut_2);
  assign _zz__29_3_inner_macOut_2 = (($signed(_zz__29_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_3_inner_activation;
    end else begin
      io_macOut = _29_3_inner_macOut;
    end
  end

  assign _zz__29_3_inner_macOut = ($signed(_zz__zz__29_3_inner_macOut) + $signed(_zz__zz__29_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_3_inner_activation <= 8'h00;
      _29_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_3_inner_activation <= io_addInput;
      end else begin
        _29_3_inner_macOut <= _zz__29_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_930 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_2_inner_macOut;
  wire       [15:0]   _zz__zz__29_2_inner_macOut_1;
  wire       [15:0]   _zz__29_2_inner_macOut_1;
  wire       [15:0]   _zz__29_2_inner_macOut_2;
  reg        [7:0]    _29_2_inner_activation;
  reg        [7:0]    _29_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_2_inner_macOut;

  assign _zz__zz__29_2_inner_macOut = ($signed(io_mulInput) * $signed(_29_2_inner_activation));
  assign _zz__zz__29_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_2_inner_macOut)) ? 16'h007f : _zz__29_2_inner_macOut_2);
  assign _zz__29_2_inner_macOut_2 = (($signed(_zz__29_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_2_inner_activation;
    end else begin
      io_macOut = _29_2_inner_macOut;
    end
  end

  assign _zz__29_2_inner_macOut = ($signed(_zz__zz__29_2_inner_macOut) + $signed(_zz__zz__29_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_2_inner_activation <= 8'h00;
      _29_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_2_inner_activation <= io_addInput;
      end else begin
        _29_2_inner_macOut <= _zz__29_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_929 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_1_inner_macOut;
  wire       [15:0]   _zz__zz__29_1_inner_macOut_1;
  wire       [15:0]   _zz__29_1_inner_macOut_1;
  wire       [15:0]   _zz__29_1_inner_macOut_2;
  reg        [7:0]    _29_1_inner_activation;
  reg        [7:0]    _29_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_1_inner_macOut;

  assign _zz__zz__29_1_inner_macOut = ($signed(io_mulInput) * $signed(_29_1_inner_activation));
  assign _zz__zz__29_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_1_inner_macOut)) ? 16'h007f : _zz__29_1_inner_macOut_2);
  assign _zz__29_1_inner_macOut_2 = (($signed(_zz__29_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_1_inner_activation;
    end else begin
      io_macOut = _29_1_inner_macOut;
    end
  end

  assign _zz__29_1_inner_macOut = ($signed(_zz__zz__29_1_inner_macOut) + $signed(_zz__zz__29_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_1_inner_activation <= 8'h00;
      _29_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_1_inner_activation <= io_addInput;
      end else begin
        _29_1_inner_macOut <= _zz__29_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_928 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__29_0_inner_macOut;
  wire       [15:0]   _zz__zz__29_0_inner_macOut_1;
  wire       [15:0]   _zz__29_0_inner_macOut_1;
  wire       [15:0]   _zz__29_0_inner_macOut_2;
  reg        [7:0]    _29_0_inner_activation;
  reg        [7:0]    _29_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__29_0_inner_macOut;

  assign _zz__zz__29_0_inner_macOut = ($signed(io_mulInput) * $signed(_29_0_inner_activation));
  assign _zz__zz__29_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__29_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__29_0_inner_macOut)) ? 16'h007f : _zz__29_0_inner_macOut_2);
  assign _zz__29_0_inner_macOut_2 = (($signed(_zz__29_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__29_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _29_0_inner_activation;
    end else begin
      io_macOut = _29_0_inner_macOut;
    end
  end

  assign _zz__29_0_inner_macOut = ($signed(_zz__zz__29_0_inner_macOut) + $signed(_zz__zz__29_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _29_0_inner_activation <= 8'h00;
      _29_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _29_0_inner_activation <= io_addInput;
      end else begin
        _29_0_inner_macOut <= _zz__29_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_927 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_31_inner_macOut;
  wire       [15:0]   _zz__zz__28_31_inner_macOut_1;
  wire       [15:0]   _zz__28_31_inner_macOut_1;
  wire       [15:0]   _zz__28_31_inner_macOut_2;
  reg        [7:0]    _28_31_inner_activation;
  reg        [7:0]    _28_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_31_inner_macOut;

  assign _zz__zz__28_31_inner_macOut = ($signed(io_mulInput) * $signed(_28_31_inner_activation));
  assign _zz__zz__28_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_31_inner_macOut)) ? 16'h007f : _zz__28_31_inner_macOut_2);
  assign _zz__28_31_inner_macOut_2 = (($signed(_zz__28_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_31_inner_activation;
    end else begin
      io_macOut = _28_31_inner_macOut;
    end
  end

  assign _zz__28_31_inner_macOut = ($signed(_zz__zz__28_31_inner_macOut) + $signed(_zz__zz__28_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_31_inner_activation <= 8'h00;
      _28_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_31_inner_activation <= io_addInput;
      end else begin
        _28_31_inner_macOut <= _zz__28_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_926 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_30_inner_macOut;
  wire       [15:0]   _zz__zz__28_30_inner_macOut_1;
  wire       [15:0]   _zz__28_30_inner_macOut_1;
  wire       [15:0]   _zz__28_30_inner_macOut_2;
  reg        [7:0]    _28_30_inner_activation;
  reg        [7:0]    _28_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_30_inner_macOut;

  assign _zz__zz__28_30_inner_macOut = ($signed(io_mulInput) * $signed(_28_30_inner_activation));
  assign _zz__zz__28_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_30_inner_macOut)) ? 16'h007f : _zz__28_30_inner_macOut_2);
  assign _zz__28_30_inner_macOut_2 = (($signed(_zz__28_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_30_inner_activation;
    end else begin
      io_macOut = _28_30_inner_macOut;
    end
  end

  assign _zz__28_30_inner_macOut = ($signed(_zz__zz__28_30_inner_macOut) + $signed(_zz__zz__28_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_30_inner_activation <= 8'h00;
      _28_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_30_inner_activation <= io_addInput;
      end else begin
        _28_30_inner_macOut <= _zz__28_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_925 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_29_inner_macOut;
  wire       [15:0]   _zz__zz__28_29_inner_macOut_1;
  wire       [15:0]   _zz__28_29_inner_macOut_1;
  wire       [15:0]   _zz__28_29_inner_macOut_2;
  reg        [7:0]    _28_29_inner_activation;
  reg        [7:0]    _28_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_29_inner_macOut;

  assign _zz__zz__28_29_inner_macOut = ($signed(io_mulInput) * $signed(_28_29_inner_activation));
  assign _zz__zz__28_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_29_inner_macOut)) ? 16'h007f : _zz__28_29_inner_macOut_2);
  assign _zz__28_29_inner_macOut_2 = (($signed(_zz__28_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_29_inner_activation;
    end else begin
      io_macOut = _28_29_inner_macOut;
    end
  end

  assign _zz__28_29_inner_macOut = ($signed(_zz__zz__28_29_inner_macOut) + $signed(_zz__zz__28_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_29_inner_activation <= 8'h00;
      _28_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_29_inner_activation <= io_addInput;
      end else begin
        _28_29_inner_macOut <= _zz__28_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_924 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_28_inner_macOut;
  wire       [15:0]   _zz__zz__28_28_inner_macOut_1;
  wire       [15:0]   _zz__28_28_inner_macOut_1;
  wire       [15:0]   _zz__28_28_inner_macOut_2;
  reg        [7:0]    _28_28_inner_activation;
  reg        [7:0]    _28_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_28_inner_macOut;

  assign _zz__zz__28_28_inner_macOut = ($signed(io_mulInput) * $signed(_28_28_inner_activation));
  assign _zz__zz__28_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_28_inner_macOut)) ? 16'h007f : _zz__28_28_inner_macOut_2);
  assign _zz__28_28_inner_macOut_2 = (($signed(_zz__28_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_28_inner_activation;
    end else begin
      io_macOut = _28_28_inner_macOut;
    end
  end

  assign _zz__28_28_inner_macOut = ($signed(_zz__zz__28_28_inner_macOut) + $signed(_zz__zz__28_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_28_inner_activation <= 8'h00;
      _28_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_28_inner_activation <= io_addInput;
      end else begin
        _28_28_inner_macOut <= _zz__28_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_923 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_27_inner_macOut;
  wire       [15:0]   _zz__zz__28_27_inner_macOut_1;
  wire       [15:0]   _zz__28_27_inner_macOut_1;
  wire       [15:0]   _zz__28_27_inner_macOut_2;
  reg        [7:0]    _28_27_inner_activation;
  reg        [7:0]    _28_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_27_inner_macOut;

  assign _zz__zz__28_27_inner_macOut = ($signed(io_mulInput) * $signed(_28_27_inner_activation));
  assign _zz__zz__28_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_27_inner_macOut)) ? 16'h007f : _zz__28_27_inner_macOut_2);
  assign _zz__28_27_inner_macOut_2 = (($signed(_zz__28_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_27_inner_activation;
    end else begin
      io_macOut = _28_27_inner_macOut;
    end
  end

  assign _zz__28_27_inner_macOut = ($signed(_zz__zz__28_27_inner_macOut) + $signed(_zz__zz__28_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_27_inner_activation <= 8'h00;
      _28_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_27_inner_activation <= io_addInput;
      end else begin
        _28_27_inner_macOut <= _zz__28_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_922 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_26_inner_macOut;
  wire       [15:0]   _zz__zz__28_26_inner_macOut_1;
  wire       [15:0]   _zz__28_26_inner_macOut_1;
  wire       [15:0]   _zz__28_26_inner_macOut_2;
  reg        [7:0]    _28_26_inner_activation;
  reg        [7:0]    _28_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_26_inner_macOut;

  assign _zz__zz__28_26_inner_macOut = ($signed(io_mulInput) * $signed(_28_26_inner_activation));
  assign _zz__zz__28_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_26_inner_macOut)) ? 16'h007f : _zz__28_26_inner_macOut_2);
  assign _zz__28_26_inner_macOut_2 = (($signed(_zz__28_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_26_inner_activation;
    end else begin
      io_macOut = _28_26_inner_macOut;
    end
  end

  assign _zz__28_26_inner_macOut = ($signed(_zz__zz__28_26_inner_macOut) + $signed(_zz__zz__28_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_26_inner_activation <= 8'h00;
      _28_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_26_inner_activation <= io_addInput;
      end else begin
        _28_26_inner_macOut <= _zz__28_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_921 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_25_inner_macOut;
  wire       [15:0]   _zz__zz__28_25_inner_macOut_1;
  wire       [15:0]   _zz__28_25_inner_macOut_1;
  wire       [15:0]   _zz__28_25_inner_macOut_2;
  reg        [7:0]    _28_25_inner_activation;
  reg        [7:0]    _28_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_25_inner_macOut;

  assign _zz__zz__28_25_inner_macOut = ($signed(io_mulInput) * $signed(_28_25_inner_activation));
  assign _zz__zz__28_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_25_inner_macOut)) ? 16'h007f : _zz__28_25_inner_macOut_2);
  assign _zz__28_25_inner_macOut_2 = (($signed(_zz__28_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_25_inner_activation;
    end else begin
      io_macOut = _28_25_inner_macOut;
    end
  end

  assign _zz__28_25_inner_macOut = ($signed(_zz__zz__28_25_inner_macOut) + $signed(_zz__zz__28_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_25_inner_activation <= 8'h00;
      _28_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_25_inner_activation <= io_addInput;
      end else begin
        _28_25_inner_macOut <= _zz__28_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_920 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_24_inner_macOut;
  wire       [15:0]   _zz__zz__28_24_inner_macOut_1;
  wire       [15:0]   _zz__28_24_inner_macOut_1;
  wire       [15:0]   _zz__28_24_inner_macOut_2;
  reg        [7:0]    _28_24_inner_activation;
  reg        [7:0]    _28_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_24_inner_macOut;

  assign _zz__zz__28_24_inner_macOut = ($signed(io_mulInput) * $signed(_28_24_inner_activation));
  assign _zz__zz__28_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_24_inner_macOut)) ? 16'h007f : _zz__28_24_inner_macOut_2);
  assign _zz__28_24_inner_macOut_2 = (($signed(_zz__28_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_24_inner_activation;
    end else begin
      io_macOut = _28_24_inner_macOut;
    end
  end

  assign _zz__28_24_inner_macOut = ($signed(_zz__zz__28_24_inner_macOut) + $signed(_zz__zz__28_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_24_inner_activation <= 8'h00;
      _28_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_24_inner_activation <= io_addInput;
      end else begin
        _28_24_inner_macOut <= _zz__28_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_919 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_23_inner_macOut;
  wire       [15:0]   _zz__zz__28_23_inner_macOut_1;
  wire       [15:0]   _zz__28_23_inner_macOut_1;
  wire       [15:0]   _zz__28_23_inner_macOut_2;
  reg        [7:0]    _28_23_inner_activation;
  reg        [7:0]    _28_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_23_inner_macOut;

  assign _zz__zz__28_23_inner_macOut = ($signed(io_mulInput) * $signed(_28_23_inner_activation));
  assign _zz__zz__28_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_23_inner_macOut)) ? 16'h007f : _zz__28_23_inner_macOut_2);
  assign _zz__28_23_inner_macOut_2 = (($signed(_zz__28_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_23_inner_activation;
    end else begin
      io_macOut = _28_23_inner_macOut;
    end
  end

  assign _zz__28_23_inner_macOut = ($signed(_zz__zz__28_23_inner_macOut) + $signed(_zz__zz__28_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_23_inner_activation <= 8'h00;
      _28_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_23_inner_activation <= io_addInput;
      end else begin
        _28_23_inner_macOut <= _zz__28_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_918 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_22_inner_macOut;
  wire       [15:0]   _zz__zz__28_22_inner_macOut_1;
  wire       [15:0]   _zz__28_22_inner_macOut_1;
  wire       [15:0]   _zz__28_22_inner_macOut_2;
  reg        [7:0]    _28_22_inner_activation;
  reg        [7:0]    _28_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_22_inner_macOut;

  assign _zz__zz__28_22_inner_macOut = ($signed(io_mulInput) * $signed(_28_22_inner_activation));
  assign _zz__zz__28_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_22_inner_macOut)) ? 16'h007f : _zz__28_22_inner_macOut_2);
  assign _zz__28_22_inner_macOut_2 = (($signed(_zz__28_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_22_inner_activation;
    end else begin
      io_macOut = _28_22_inner_macOut;
    end
  end

  assign _zz__28_22_inner_macOut = ($signed(_zz__zz__28_22_inner_macOut) + $signed(_zz__zz__28_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_22_inner_activation <= 8'h00;
      _28_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_22_inner_activation <= io_addInput;
      end else begin
        _28_22_inner_macOut <= _zz__28_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_917 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_21_inner_macOut;
  wire       [15:0]   _zz__zz__28_21_inner_macOut_1;
  wire       [15:0]   _zz__28_21_inner_macOut_1;
  wire       [15:0]   _zz__28_21_inner_macOut_2;
  reg        [7:0]    _28_21_inner_activation;
  reg        [7:0]    _28_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_21_inner_macOut;

  assign _zz__zz__28_21_inner_macOut = ($signed(io_mulInput) * $signed(_28_21_inner_activation));
  assign _zz__zz__28_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_21_inner_macOut)) ? 16'h007f : _zz__28_21_inner_macOut_2);
  assign _zz__28_21_inner_macOut_2 = (($signed(_zz__28_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_21_inner_activation;
    end else begin
      io_macOut = _28_21_inner_macOut;
    end
  end

  assign _zz__28_21_inner_macOut = ($signed(_zz__zz__28_21_inner_macOut) + $signed(_zz__zz__28_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_21_inner_activation <= 8'h00;
      _28_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_21_inner_activation <= io_addInput;
      end else begin
        _28_21_inner_macOut <= _zz__28_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_916 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_20_inner_macOut;
  wire       [15:0]   _zz__zz__28_20_inner_macOut_1;
  wire       [15:0]   _zz__28_20_inner_macOut_1;
  wire       [15:0]   _zz__28_20_inner_macOut_2;
  reg        [7:0]    _28_20_inner_activation;
  reg        [7:0]    _28_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_20_inner_macOut;

  assign _zz__zz__28_20_inner_macOut = ($signed(io_mulInput) * $signed(_28_20_inner_activation));
  assign _zz__zz__28_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_20_inner_macOut)) ? 16'h007f : _zz__28_20_inner_macOut_2);
  assign _zz__28_20_inner_macOut_2 = (($signed(_zz__28_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_20_inner_activation;
    end else begin
      io_macOut = _28_20_inner_macOut;
    end
  end

  assign _zz__28_20_inner_macOut = ($signed(_zz__zz__28_20_inner_macOut) + $signed(_zz__zz__28_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_20_inner_activation <= 8'h00;
      _28_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_20_inner_activation <= io_addInput;
      end else begin
        _28_20_inner_macOut <= _zz__28_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_915 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_19_inner_macOut;
  wire       [15:0]   _zz__zz__28_19_inner_macOut_1;
  wire       [15:0]   _zz__28_19_inner_macOut_1;
  wire       [15:0]   _zz__28_19_inner_macOut_2;
  reg        [7:0]    _28_19_inner_activation;
  reg        [7:0]    _28_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_19_inner_macOut;

  assign _zz__zz__28_19_inner_macOut = ($signed(io_mulInput) * $signed(_28_19_inner_activation));
  assign _zz__zz__28_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_19_inner_macOut)) ? 16'h007f : _zz__28_19_inner_macOut_2);
  assign _zz__28_19_inner_macOut_2 = (($signed(_zz__28_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_19_inner_activation;
    end else begin
      io_macOut = _28_19_inner_macOut;
    end
  end

  assign _zz__28_19_inner_macOut = ($signed(_zz__zz__28_19_inner_macOut) + $signed(_zz__zz__28_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_19_inner_activation <= 8'h00;
      _28_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_19_inner_activation <= io_addInput;
      end else begin
        _28_19_inner_macOut <= _zz__28_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_914 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_18_inner_macOut;
  wire       [15:0]   _zz__zz__28_18_inner_macOut_1;
  wire       [15:0]   _zz__28_18_inner_macOut_1;
  wire       [15:0]   _zz__28_18_inner_macOut_2;
  reg        [7:0]    _28_18_inner_activation;
  reg        [7:0]    _28_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_18_inner_macOut;

  assign _zz__zz__28_18_inner_macOut = ($signed(io_mulInput) * $signed(_28_18_inner_activation));
  assign _zz__zz__28_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_18_inner_macOut)) ? 16'h007f : _zz__28_18_inner_macOut_2);
  assign _zz__28_18_inner_macOut_2 = (($signed(_zz__28_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_18_inner_activation;
    end else begin
      io_macOut = _28_18_inner_macOut;
    end
  end

  assign _zz__28_18_inner_macOut = ($signed(_zz__zz__28_18_inner_macOut) + $signed(_zz__zz__28_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_18_inner_activation <= 8'h00;
      _28_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_18_inner_activation <= io_addInput;
      end else begin
        _28_18_inner_macOut <= _zz__28_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_913 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_17_inner_macOut;
  wire       [15:0]   _zz__zz__28_17_inner_macOut_1;
  wire       [15:0]   _zz__28_17_inner_macOut_1;
  wire       [15:0]   _zz__28_17_inner_macOut_2;
  reg        [7:0]    _28_17_inner_activation;
  reg        [7:0]    _28_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_17_inner_macOut;

  assign _zz__zz__28_17_inner_macOut = ($signed(io_mulInput) * $signed(_28_17_inner_activation));
  assign _zz__zz__28_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_17_inner_macOut)) ? 16'h007f : _zz__28_17_inner_macOut_2);
  assign _zz__28_17_inner_macOut_2 = (($signed(_zz__28_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_17_inner_activation;
    end else begin
      io_macOut = _28_17_inner_macOut;
    end
  end

  assign _zz__28_17_inner_macOut = ($signed(_zz__zz__28_17_inner_macOut) + $signed(_zz__zz__28_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_17_inner_activation <= 8'h00;
      _28_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_17_inner_activation <= io_addInput;
      end else begin
        _28_17_inner_macOut <= _zz__28_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_912 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_16_inner_macOut;
  wire       [15:0]   _zz__zz__28_16_inner_macOut_1;
  wire       [15:0]   _zz__28_16_inner_macOut_1;
  wire       [15:0]   _zz__28_16_inner_macOut_2;
  reg        [7:0]    _28_16_inner_activation;
  reg        [7:0]    _28_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_16_inner_macOut;

  assign _zz__zz__28_16_inner_macOut = ($signed(io_mulInput) * $signed(_28_16_inner_activation));
  assign _zz__zz__28_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_16_inner_macOut)) ? 16'h007f : _zz__28_16_inner_macOut_2);
  assign _zz__28_16_inner_macOut_2 = (($signed(_zz__28_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_16_inner_activation;
    end else begin
      io_macOut = _28_16_inner_macOut;
    end
  end

  assign _zz__28_16_inner_macOut = ($signed(_zz__zz__28_16_inner_macOut) + $signed(_zz__zz__28_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_16_inner_activation <= 8'h00;
      _28_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_16_inner_activation <= io_addInput;
      end else begin
        _28_16_inner_macOut <= _zz__28_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_911 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_15_inner_macOut;
  wire       [15:0]   _zz__zz__28_15_inner_macOut_1;
  wire       [15:0]   _zz__28_15_inner_macOut_1;
  wire       [15:0]   _zz__28_15_inner_macOut_2;
  reg        [7:0]    _28_15_inner_activation;
  reg        [7:0]    _28_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_15_inner_macOut;

  assign _zz__zz__28_15_inner_macOut = ($signed(io_mulInput) * $signed(_28_15_inner_activation));
  assign _zz__zz__28_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_15_inner_macOut)) ? 16'h007f : _zz__28_15_inner_macOut_2);
  assign _zz__28_15_inner_macOut_2 = (($signed(_zz__28_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_15_inner_activation;
    end else begin
      io_macOut = _28_15_inner_macOut;
    end
  end

  assign _zz__28_15_inner_macOut = ($signed(_zz__zz__28_15_inner_macOut) + $signed(_zz__zz__28_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_15_inner_activation <= 8'h00;
      _28_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_15_inner_activation <= io_addInput;
      end else begin
        _28_15_inner_macOut <= _zz__28_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_910 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_14_inner_macOut;
  wire       [15:0]   _zz__zz__28_14_inner_macOut_1;
  wire       [15:0]   _zz__28_14_inner_macOut_1;
  wire       [15:0]   _zz__28_14_inner_macOut_2;
  reg        [7:0]    _28_14_inner_activation;
  reg        [7:0]    _28_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_14_inner_macOut;

  assign _zz__zz__28_14_inner_macOut = ($signed(io_mulInput) * $signed(_28_14_inner_activation));
  assign _zz__zz__28_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_14_inner_macOut)) ? 16'h007f : _zz__28_14_inner_macOut_2);
  assign _zz__28_14_inner_macOut_2 = (($signed(_zz__28_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_14_inner_activation;
    end else begin
      io_macOut = _28_14_inner_macOut;
    end
  end

  assign _zz__28_14_inner_macOut = ($signed(_zz__zz__28_14_inner_macOut) + $signed(_zz__zz__28_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_14_inner_activation <= 8'h00;
      _28_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_14_inner_activation <= io_addInput;
      end else begin
        _28_14_inner_macOut <= _zz__28_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_909 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_13_inner_macOut;
  wire       [15:0]   _zz__zz__28_13_inner_macOut_1;
  wire       [15:0]   _zz__28_13_inner_macOut_1;
  wire       [15:0]   _zz__28_13_inner_macOut_2;
  reg        [7:0]    _28_13_inner_activation;
  reg        [7:0]    _28_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_13_inner_macOut;

  assign _zz__zz__28_13_inner_macOut = ($signed(io_mulInput) * $signed(_28_13_inner_activation));
  assign _zz__zz__28_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_13_inner_macOut)) ? 16'h007f : _zz__28_13_inner_macOut_2);
  assign _zz__28_13_inner_macOut_2 = (($signed(_zz__28_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_13_inner_activation;
    end else begin
      io_macOut = _28_13_inner_macOut;
    end
  end

  assign _zz__28_13_inner_macOut = ($signed(_zz__zz__28_13_inner_macOut) + $signed(_zz__zz__28_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_13_inner_activation <= 8'h00;
      _28_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_13_inner_activation <= io_addInput;
      end else begin
        _28_13_inner_macOut <= _zz__28_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_908 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_12_inner_macOut;
  wire       [15:0]   _zz__zz__28_12_inner_macOut_1;
  wire       [15:0]   _zz__28_12_inner_macOut_1;
  wire       [15:0]   _zz__28_12_inner_macOut_2;
  reg        [7:0]    _28_12_inner_activation;
  reg        [7:0]    _28_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_12_inner_macOut;

  assign _zz__zz__28_12_inner_macOut = ($signed(io_mulInput) * $signed(_28_12_inner_activation));
  assign _zz__zz__28_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_12_inner_macOut)) ? 16'h007f : _zz__28_12_inner_macOut_2);
  assign _zz__28_12_inner_macOut_2 = (($signed(_zz__28_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_12_inner_activation;
    end else begin
      io_macOut = _28_12_inner_macOut;
    end
  end

  assign _zz__28_12_inner_macOut = ($signed(_zz__zz__28_12_inner_macOut) + $signed(_zz__zz__28_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_12_inner_activation <= 8'h00;
      _28_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_12_inner_activation <= io_addInput;
      end else begin
        _28_12_inner_macOut <= _zz__28_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_907 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_11_inner_macOut;
  wire       [15:0]   _zz__zz__28_11_inner_macOut_1;
  wire       [15:0]   _zz__28_11_inner_macOut_1;
  wire       [15:0]   _zz__28_11_inner_macOut_2;
  reg        [7:0]    _28_11_inner_activation;
  reg        [7:0]    _28_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_11_inner_macOut;

  assign _zz__zz__28_11_inner_macOut = ($signed(io_mulInput) * $signed(_28_11_inner_activation));
  assign _zz__zz__28_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_11_inner_macOut)) ? 16'h007f : _zz__28_11_inner_macOut_2);
  assign _zz__28_11_inner_macOut_2 = (($signed(_zz__28_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_11_inner_activation;
    end else begin
      io_macOut = _28_11_inner_macOut;
    end
  end

  assign _zz__28_11_inner_macOut = ($signed(_zz__zz__28_11_inner_macOut) + $signed(_zz__zz__28_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_11_inner_activation <= 8'h00;
      _28_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_11_inner_activation <= io_addInput;
      end else begin
        _28_11_inner_macOut <= _zz__28_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_906 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_10_inner_macOut;
  wire       [15:0]   _zz__zz__28_10_inner_macOut_1;
  wire       [15:0]   _zz__28_10_inner_macOut_1;
  wire       [15:0]   _zz__28_10_inner_macOut_2;
  reg        [7:0]    _28_10_inner_activation;
  reg        [7:0]    _28_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_10_inner_macOut;

  assign _zz__zz__28_10_inner_macOut = ($signed(io_mulInput) * $signed(_28_10_inner_activation));
  assign _zz__zz__28_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_10_inner_macOut)) ? 16'h007f : _zz__28_10_inner_macOut_2);
  assign _zz__28_10_inner_macOut_2 = (($signed(_zz__28_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_10_inner_activation;
    end else begin
      io_macOut = _28_10_inner_macOut;
    end
  end

  assign _zz__28_10_inner_macOut = ($signed(_zz__zz__28_10_inner_macOut) + $signed(_zz__zz__28_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_10_inner_activation <= 8'h00;
      _28_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_10_inner_activation <= io_addInput;
      end else begin
        _28_10_inner_macOut <= _zz__28_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_905 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_9_inner_macOut;
  wire       [15:0]   _zz__zz__28_9_inner_macOut_1;
  wire       [15:0]   _zz__28_9_inner_macOut_1;
  wire       [15:0]   _zz__28_9_inner_macOut_2;
  reg        [7:0]    _28_9_inner_activation;
  reg        [7:0]    _28_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_9_inner_macOut;

  assign _zz__zz__28_9_inner_macOut = ($signed(io_mulInput) * $signed(_28_9_inner_activation));
  assign _zz__zz__28_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_9_inner_macOut)) ? 16'h007f : _zz__28_9_inner_macOut_2);
  assign _zz__28_9_inner_macOut_2 = (($signed(_zz__28_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_9_inner_activation;
    end else begin
      io_macOut = _28_9_inner_macOut;
    end
  end

  assign _zz__28_9_inner_macOut = ($signed(_zz__zz__28_9_inner_macOut) + $signed(_zz__zz__28_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_9_inner_activation <= 8'h00;
      _28_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_9_inner_activation <= io_addInput;
      end else begin
        _28_9_inner_macOut <= _zz__28_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_904 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_8_inner_macOut;
  wire       [15:0]   _zz__zz__28_8_inner_macOut_1;
  wire       [15:0]   _zz__28_8_inner_macOut_1;
  wire       [15:0]   _zz__28_8_inner_macOut_2;
  reg        [7:0]    _28_8_inner_activation;
  reg        [7:0]    _28_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_8_inner_macOut;

  assign _zz__zz__28_8_inner_macOut = ($signed(io_mulInput) * $signed(_28_8_inner_activation));
  assign _zz__zz__28_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_8_inner_macOut)) ? 16'h007f : _zz__28_8_inner_macOut_2);
  assign _zz__28_8_inner_macOut_2 = (($signed(_zz__28_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_8_inner_activation;
    end else begin
      io_macOut = _28_8_inner_macOut;
    end
  end

  assign _zz__28_8_inner_macOut = ($signed(_zz__zz__28_8_inner_macOut) + $signed(_zz__zz__28_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_8_inner_activation <= 8'h00;
      _28_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_8_inner_activation <= io_addInput;
      end else begin
        _28_8_inner_macOut <= _zz__28_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_903 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_7_inner_macOut;
  wire       [15:0]   _zz__zz__28_7_inner_macOut_1;
  wire       [15:0]   _zz__28_7_inner_macOut_1;
  wire       [15:0]   _zz__28_7_inner_macOut_2;
  reg        [7:0]    _28_7_inner_activation;
  reg        [7:0]    _28_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_7_inner_macOut;

  assign _zz__zz__28_7_inner_macOut = ($signed(io_mulInput) * $signed(_28_7_inner_activation));
  assign _zz__zz__28_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_7_inner_macOut)) ? 16'h007f : _zz__28_7_inner_macOut_2);
  assign _zz__28_7_inner_macOut_2 = (($signed(_zz__28_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_7_inner_activation;
    end else begin
      io_macOut = _28_7_inner_macOut;
    end
  end

  assign _zz__28_7_inner_macOut = ($signed(_zz__zz__28_7_inner_macOut) + $signed(_zz__zz__28_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_7_inner_activation <= 8'h00;
      _28_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_7_inner_activation <= io_addInput;
      end else begin
        _28_7_inner_macOut <= _zz__28_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_902 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_6_inner_macOut;
  wire       [15:0]   _zz__zz__28_6_inner_macOut_1;
  wire       [15:0]   _zz__28_6_inner_macOut_1;
  wire       [15:0]   _zz__28_6_inner_macOut_2;
  reg        [7:0]    _28_6_inner_activation;
  reg        [7:0]    _28_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_6_inner_macOut;

  assign _zz__zz__28_6_inner_macOut = ($signed(io_mulInput) * $signed(_28_6_inner_activation));
  assign _zz__zz__28_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_6_inner_macOut)) ? 16'h007f : _zz__28_6_inner_macOut_2);
  assign _zz__28_6_inner_macOut_2 = (($signed(_zz__28_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_6_inner_activation;
    end else begin
      io_macOut = _28_6_inner_macOut;
    end
  end

  assign _zz__28_6_inner_macOut = ($signed(_zz__zz__28_6_inner_macOut) + $signed(_zz__zz__28_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_6_inner_activation <= 8'h00;
      _28_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_6_inner_activation <= io_addInput;
      end else begin
        _28_6_inner_macOut <= _zz__28_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_901 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_5_inner_macOut;
  wire       [15:0]   _zz__zz__28_5_inner_macOut_1;
  wire       [15:0]   _zz__28_5_inner_macOut_1;
  wire       [15:0]   _zz__28_5_inner_macOut_2;
  reg        [7:0]    _28_5_inner_activation;
  reg        [7:0]    _28_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_5_inner_macOut;

  assign _zz__zz__28_5_inner_macOut = ($signed(io_mulInput) * $signed(_28_5_inner_activation));
  assign _zz__zz__28_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_5_inner_macOut)) ? 16'h007f : _zz__28_5_inner_macOut_2);
  assign _zz__28_5_inner_macOut_2 = (($signed(_zz__28_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_5_inner_activation;
    end else begin
      io_macOut = _28_5_inner_macOut;
    end
  end

  assign _zz__28_5_inner_macOut = ($signed(_zz__zz__28_5_inner_macOut) + $signed(_zz__zz__28_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_5_inner_activation <= 8'h00;
      _28_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_5_inner_activation <= io_addInput;
      end else begin
        _28_5_inner_macOut <= _zz__28_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_900 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_4_inner_macOut;
  wire       [15:0]   _zz__zz__28_4_inner_macOut_1;
  wire       [15:0]   _zz__28_4_inner_macOut_1;
  wire       [15:0]   _zz__28_4_inner_macOut_2;
  reg        [7:0]    _28_4_inner_activation;
  reg        [7:0]    _28_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_4_inner_macOut;

  assign _zz__zz__28_4_inner_macOut = ($signed(io_mulInput) * $signed(_28_4_inner_activation));
  assign _zz__zz__28_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_4_inner_macOut)) ? 16'h007f : _zz__28_4_inner_macOut_2);
  assign _zz__28_4_inner_macOut_2 = (($signed(_zz__28_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_4_inner_activation;
    end else begin
      io_macOut = _28_4_inner_macOut;
    end
  end

  assign _zz__28_4_inner_macOut = ($signed(_zz__zz__28_4_inner_macOut) + $signed(_zz__zz__28_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_4_inner_activation <= 8'h00;
      _28_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_4_inner_activation <= io_addInput;
      end else begin
        _28_4_inner_macOut <= _zz__28_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_899 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_3_inner_macOut;
  wire       [15:0]   _zz__zz__28_3_inner_macOut_1;
  wire       [15:0]   _zz__28_3_inner_macOut_1;
  wire       [15:0]   _zz__28_3_inner_macOut_2;
  reg        [7:0]    _28_3_inner_activation;
  reg        [7:0]    _28_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_3_inner_macOut;

  assign _zz__zz__28_3_inner_macOut = ($signed(io_mulInput) * $signed(_28_3_inner_activation));
  assign _zz__zz__28_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_3_inner_macOut)) ? 16'h007f : _zz__28_3_inner_macOut_2);
  assign _zz__28_3_inner_macOut_2 = (($signed(_zz__28_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_3_inner_activation;
    end else begin
      io_macOut = _28_3_inner_macOut;
    end
  end

  assign _zz__28_3_inner_macOut = ($signed(_zz__zz__28_3_inner_macOut) + $signed(_zz__zz__28_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_3_inner_activation <= 8'h00;
      _28_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_3_inner_activation <= io_addInput;
      end else begin
        _28_3_inner_macOut <= _zz__28_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_898 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_2_inner_macOut;
  wire       [15:0]   _zz__zz__28_2_inner_macOut_1;
  wire       [15:0]   _zz__28_2_inner_macOut_1;
  wire       [15:0]   _zz__28_2_inner_macOut_2;
  reg        [7:0]    _28_2_inner_activation;
  reg        [7:0]    _28_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_2_inner_macOut;

  assign _zz__zz__28_2_inner_macOut = ($signed(io_mulInput) * $signed(_28_2_inner_activation));
  assign _zz__zz__28_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_2_inner_macOut)) ? 16'h007f : _zz__28_2_inner_macOut_2);
  assign _zz__28_2_inner_macOut_2 = (($signed(_zz__28_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_2_inner_activation;
    end else begin
      io_macOut = _28_2_inner_macOut;
    end
  end

  assign _zz__28_2_inner_macOut = ($signed(_zz__zz__28_2_inner_macOut) + $signed(_zz__zz__28_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_2_inner_activation <= 8'h00;
      _28_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_2_inner_activation <= io_addInput;
      end else begin
        _28_2_inner_macOut <= _zz__28_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_897 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_1_inner_macOut;
  wire       [15:0]   _zz__zz__28_1_inner_macOut_1;
  wire       [15:0]   _zz__28_1_inner_macOut_1;
  wire       [15:0]   _zz__28_1_inner_macOut_2;
  reg        [7:0]    _28_1_inner_activation;
  reg        [7:0]    _28_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_1_inner_macOut;

  assign _zz__zz__28_1_inner_macOut = ($signed(io_mulInput) * $signed(_28_1_inner_activation));
  assign _zz__zz__28_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_1_inner_macOut)) ? 16'h007f : _zz__28_1_inner_macOut_2);
  assign _zz__28_1_inner_macOut_2 = (($signed(_zz__28_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_1_inner_activation;
    end else begin
      io_macOut = _28_1_inner_macOut;
    end
  end

  assign _zz__28_1_inner_macOut = ($signed(_zz__zz__28_1_inner_macOut) + $signed(_zz__zz__28_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_1_inner_activation <= 8'h00;
      _28_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_1_inner_activation <= io_addInput;
      end else begin
        _28_1_inner_macOut <= _zz__28_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_896 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__28_0_inner_macOut;
  wire       [15:0]   _zz__zz__28_0_inner_macOut_1;
  wire       [15:0]   _zz__28_0_inner_macOut_1;
  wire       [15:0]   _zz__28_0_inner_macOut_2;
  reg        [7:0]    _28_0_inner_activation;
  reg        [7:0]    _28_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__28_0_inner_macOut;

  assign _zz__zz__28_0_inner_macOut = ($signed(io_mulInput) * $signed(_28_0_inner_activation));
  assign _zz__zz__28_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__28_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__28_0_inner_macOut)) ? 16'h007f : _zz__28_0_inner_macOut_2);
  assign _zz__28_0_inner_macOut_2 = (($signed(_zz__28_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__28_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _28_0_inner_activation;
    end else begin
      io_macOut = _28_0_inner_macOut;
    end
  end

  assign _zz__28_0_inner_macOut = ($signed(_zz__zz__28_0_inner_macOut) + $signed(_zz__zz__28_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _28_0_inner_activation <= 8'h00;
      _28_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _28_0_inner_activation <= io_addInput;
      end else begin
        _28_0_inner_macOut <= _zz__28_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_895 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_31_inner_macOut;
  wire       [15:0]   _zz__zz__27_31_inner_macOut_1;
  wire       [15:0]   _zz__27_31_inner_macOut_1;
  wire       [15:0]   _zz__27_31_inner_macOut_2;
  reg        [7:0]    _27_31_inner_activation;
  reg        [7:0]    _27_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_31_inner_macOut;

  assign _zz__zz__27_31_inner_macOut = ($signed(io_mulInput) * $signed(_27_31_inner_activation));
  assign _zz__zz__27_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_31_inner_macOut)) ? 16'h007f : _zz__27_31_inner_macOut_2);
  assign _zz__27_31_inner_macOut_2 = (($signed(_zz__27_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_31_inner_activation;
    end else begin
      io_macOut = _27_31_inner_macOut;
    end
  end

  assign _zz__27_31_inner_macOut = ($signed(_zz__zz__27_31_inner_macOut) + $signed(_zz__zz__27_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_31_inner_activation <= 8'h00;
      _27_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_31_inner_activation <= io_addInput;
      end else begin
        _27_31_inner_macOut <= _zz__27_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_894 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_30_inner_macOut;
  wire       [15:0]   _zz__zz__27_30_inner_macOut_1;
  wire       [15:0]   _zz__27_30_inner_macOut_1;
  wire       [15:0]   _zz__27_30_inner_macOut_2;
  reg        [7:0]    _27_30_inner_activation;
  reg        [7:0]    _27_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_30_inner_macOut;

  assign _zz__zz__27_30_inner_macOut = ($signed(io_mulInput) * $signed(_27_30_inner_activation));
  assign _zz__zz__27_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_30_inner_macOut)) ? 16'h007f : _zz__27_30_inner_macOut_2);
  assign _zz__27_30_inner_macOut_2 = (($signed(_zz__27_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_30_inner_activation;
    end else begin
      io_macOut = _27_30_inner_macOut;
    end
  end

  assign _zz__27_30_inner_macOut = ($signed(_zz__zz__27_30_inner_macOut) + $signed(_zz__zz__27_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_30_inner_activation <= 8'h00;
      _27_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_30_inner_activation <= io_addInput;
      end else begin
        _27_30_inner_macOut <= _zz__27_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_893 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_29_inner_macOut;
  wire       [15:0]   _zz__zz__27_29_inner_macOut_1;
  wire       [15:0]   _zz__27_29_inner_macOut_1;
  wire       [15:0]   _zz__27_29_inner_macOut_2;
  reg        [7:0]    _27_29_inner_activation;
  reg        [7:0]    _27_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_29_inner_macOut;

  assign _zz__zz__27_29_inner_macOut = ($signed(io_mulInput) * $signed(_27_29_inner_activation));
  assign _zz__zz__27_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_29_inner_macOut)) ? 16'h007f : _zz__27_29_inner_macOut_2);
  assign _zz__27_29_inner_macOut_2 = (($signed(_zz__27_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_29_inner_activation;
    end else begin
      io_macOut = _27_29_inner_macOut;
    end
  end

  assign _zz__27_29_inner_macOut = ($signed(_zz__zz__27_29_inner_macOut) + $signed(_zz__zz__27_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_29_inner_activation <= 8'h00;
      _27_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_29_inner_activation <= io_addInput;
      end else begin
        _27_29_inner_macOut <= _zz__27_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_892 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_28_inner_macOut;
  wire       [15:0]   _zz__zz__27_28_inner_macOut_1;
  wire       [15:0]   _zz__27_28_inner_macOut_1;
  wire       [15:0]   _zz__27_28_inner_macOut_2;
  reg        [7:0]    _27_28_inner_activation;
  reg        [7:0]    _27_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_28_inner_macOut;

  assign _zz__zz__27_28_inner_macOut = ($signed(io_mulInput) * $signed(_27_28_inner_activation));
  assign _zz__zz__27_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_28_inner_macOut)) ? 16'h007f : _zz__27_28_inner_macOut_2);
  assign _zz__27_28_inner_macOut_2 = (($signed(_zz__27_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_28_inner_activation;
    end else begin
      io_macOut = _27_28_inner_macOut;
    end
  end

  assign _zz__27_28_inner_macOut = ($signed(_zz__zz__27_28_inner_macOut) + $signed(_zz__zz__27_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_28_inner_activation <= 8'h00;
      _27_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_28_inner_activation <= io_addInput;
      end else begin
        _27_28_inner_macOut <= _zz__27_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_891 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_27_inner_macOut;
  wire       [15:0]   _zz__zz__27_27_inner_macOut_1;
  wire       [15:0]   _zz__27_27_inner_macOut_1;
  wire       [15:0]   _zz__27_27_inner_macOut_2;
  reg        [7:0]    _27_27_inner_activation;
  reg        [7:0]    _27_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_27_inner_macOut;

  assign _zz__zz__27_27_inner_macOut = ($signed(io_mulInput) * $signed(_27_27_inner_activation));
  assign _zz__zz__27_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_27_inner_macOut)) ? 16'h007f : _zz__27_27_inner_macOut_2);
  assign _zz__27_27_inner_macOut_2 = (($signed(_zz__27_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_27_inner_activation;
    end else begin
      io_macOut = _27_27_inner_macOut;
    end
  end

  assign _zz__27_27_inner_macOut = ($signed(_zz__zz__27_27_inner_macOut) + $signed(_zz__zz__27_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_27_inner_activation <= 8'h00;
      _27_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_27_inner_activation <= io_addInput;
      end else begin
        _27_27_inner_macOut <= _zz__27_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_890 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_26_inner_macOut;
  wire       [15:0]   _zz__zz__27_26_inner_macOut_1;
  wire       [15:0]   _zz__27_26_inner_macOut_1;
  wire       [15:0]   _zz__27_26_inner_macOut_2;
  reg        [7:0]    _27_26_inner_activation;
  reg        [7:0]    _27_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_26_inner_macOut;

  assign _zz__zz__27_26_inner_macOut = ($signed(io_mulInput) * $signed(_27_26_inner_activation));
  assign _zz__zz__27_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_26_inner_macOut)) ? 16'h007f : _zz__27_26_inner_macOut_2);
  assign _zz__27_26_inner_macOut_2 = (($signed(_zz__27_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_26_inner_activation;
    end else begin
      io_macOut = _27_26_inner_macOut;
    end
  end

  assign _zz__27_26_inner_macOut = ($signed(_zz__zz__27_26_inner_macOut) + $signed(_zz__zz__27_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_26_inner_activation <= 8'h00;
      _27_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_26_inner_activation <= io_addInput;
      end else begin
        _27_26_inner_macOut <= _zz__27_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_889 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_25_inner_macOut;
  wire       [15:0]   _zz__zz__27_25_inner_macOut_1;
  wire       [15:0]   _zz__27_25_inner_macOut_1;
  wire       [15:0]   _zz__27_25_inner_macOut_2;
  reg        [7:0]    _27_25_inner_activation;
  reg        [7:0]    _27_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_25_inner_macOut;

  assign _zz__zz__27_25_inner_macOut = ($signed(io_mulInput) * $signed(_27_25_inner_activation));
  assign _zz__zz__27_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_25_inner_macOut)) ? 16'h007f : _zz__27_25_inner_macOut_2);
  assign _zz__27_25_inner_macOut_2 = (($signed(_zz__27_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_25_inner_activation;
    end else begin
      io_macOut = _27_25_inner_macOut;
    end
  end

  assign _zz__27_25_inner_macOut = ($signed(_zz__zz__27_25_inner_macOut) + $signed(_zz__zz__27_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_25_inner_activation <= 8'h00;
      _27_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_25_inner_activation <= io_addInput;
      end else begin
        _27_25_inner_macOut <= _zz__27_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_888 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_24_inner_macOut;
  wire       [15:0]   _zz__zz__27_24_inner_macOut_1;
  wire       [15:0]   _zz__27_24_inner_macOut_1;
  wire       [15:0]   _zz__27_24_inner_macOut_2;
  reg        [7:0]    _27_24_inner_activation;
  reg        [7:0]    _27_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_24_inner_macOut;

  assign _zz__zz__27_24_inner_macOut = ($signed(io_mulInput) * $signed(_27_24_inner_activation));
  assign _zz__zz__27_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_24_inner_macOut)) ? 16'h007f : _zz__27_24_inner_macOut_2);
  assign _zz__27_24_inner_macOut_2 = (($signed(_zz__27_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_24_inner_activation;
    end else begin
      io_macOut = _27_24_inner_macOut;
    end
  end

  assign _zz__27_24_inner_macOut = ($signed(_zz__zz__27_24_inner_macOut) + $signed(_zz__zz__27_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_24_inner_activation <= 8'h00;
      _27_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_24_inner_activation <= io_addInput;
      end else begin
        _27_24_inner_macOut <= _zz__27_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_887 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_23_inner_macOut;
  wire       [15:0]   _zz__zz__27_23_inner_macOut_1;
  wire       [15:0]   _zz__27_23_inner_macOut_1;
  wire       [15:0]   _zz__27_23_inner_macOut_2;
  reg        [7:0]    _27_23_inner_activation;
  reg        [7:0]    _27_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_23_inner_macOut;

  assign _zz__zz__27_23_inner_macOut = ($signed(io_mulInput) * $signed(_27_23_inner_activation));
  assign _zz__zz__27_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_23_inner_macOut)) ? 16'h007f : _zz__27_23_inner_macOut_2);
  assign _zz__27_23_inner_macOut_2 = (($signed(_zz__27_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_23_inner_activation;
    end else begin
      io_macOut = _27_23_inner_macOut;
    end
  end

  assign _zz__27_23_inner_macOut = ($signed(_zz__zz__27_23_inner_macOut) + $signed(_zz__zz__27_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_23_inner_activation <= 8'h00;
      _27_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_23_inner_activation <= io_addInput;
      end else begin
        _27_23_inner_macOut <= _zz__27_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_886 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_22_inner_macOut;
  wire       [15:0]   _zz__zz__27_22_inner_macOut_1;
  wire       [15:0]   _zz__27_22_inner_macOut_1;
  wire       [15:0]   _zz__27_22_inner_macOut_2;
  reg        [7:0]    _27_22_inner_activation;
  reg        [7:0]    _27_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_22_inner_macOut;

  assign _zz__zz__27_22_inner_macOut = ($signed(io_mulInput) * $signed(_27_22_inner_activation));
  assign _zz__zz__27_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_22_inner_macOut)) ? 16'h007f : _zz__27_22_inner_macOut_2);
  assign _zz__27_22_inner_macOut_2 = (($signed(_zz__27_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_22_inner_activation;
    end else begin
      io_macOut = _27_22_inner_macOut;
    end
  end

  assign _zz__27_22_inner_macOut = ($signed(_zz__zz__27_22_inner_macOut) + $signed(_zz__zz__27_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_22_inner_activation <= 8'h00;
      _27_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_22_inner_activation <= io_addInput;
      end else begin
        _27_22_inner_macOut <= _zz__27_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_885 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_21_inner_macOut;
  wire       [15:0]   _zz__zz__27_21_inner_macOut_1;
  wire       [15:0]   _zz__27_21_inner_macOut_1;
  wire       [15:0]   _zz__27_21_inner_macOut_2;
  reg        [7:0]    _27_21_inner_activation;
  reg        [7:0]    _27_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_21_inner_macOut;

  assign _zz__zz__27_21_inner_macOut = ($signed(io_mulInput) * $signed(_27_21_inner_activation));
  assign _zz__zz__27_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_21_inner_macOut)) ? 16'h007f : _zz__27_21_inner_macOut_2);
  assign _zz__27_21_inner_macOut_2 = (($signed(_zz__27_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_21_inner_activation;
    end else begin
      io_macOut = _27_21_inner_macOut;
    end
  end

  assign _zz__27_21_inner_macOut = ($signed(_zz__zz__27_21_inner_macOut) + $signed(_zz__zz__27_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_21_inner_activation <= 8'h00;
      _27_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_21_inner_activation <= io_addInput;
      end else begin
        _27_21_inner_macOut <= _zz__27_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_884 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_20_inner_macOut;
  wire       [15:0]   _zz__zz__27_20_inner_macOut_1;
  wire       [15:0]   _zz__27_20_inner_macOut_1;
  wire       [15:0]   _zz__27_20_inner_macOut_2;
  reg        [7:0]    _27_20_inner_activation;
  reg        [7:0]    _27_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_20_inner_macOut;

  assign _zz__zz__27_20_inner_macOut = ($signed(io_mulInput) * $signed(_27_20_inner_activation));
  assign _zz__zz__27_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_20_inner_macOut)) ? 16'h007f : _zz__27_20_inner_macOut_2);
  assign _zz__27_20_inner_macOut_2 = (($signed(_zz__27_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_20_inner_activation;
    end else begin
      io_macOut = _27_20_inner_macOut;
    end
  end

  assign _zz__27_20_inner_macOut = ($signed(_zz__zz__27_20_inner_macOut) + $signed(_zz__zz__27_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_20_inner_activation <= 8'h00;
      _27_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_20_inner_activation <= io_addInput;
      end else begin
        _27_20_inner_macOut <= _zz__27_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_883 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_19_inner_macOut;
  wire       [15:0]   _zz__zz__27_19_inner_macOut_1;
  wire       [15:0]   _zz__27_19_inner_macOut_1;
  wire       [15:0]   _zz__27_19_inner_macOut_2;
  reg        [7:0]    _27_19_inner_activation;
  reg        [7:0]    _27_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_19_inner_macOut;

  assign _zz__zz__27_19_inner_macOut = ($signed(io_mulInput) * $signed(_27_19_inner_activation));
  assign _zz__zz__27_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_19_inner_macOut)) ? 16'h007f : _zz__27_19_inner_macOut_2);
  assign _zz__27_19_inner_macOut_2 = (($signed(_zz__27_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_19_inner_activation;
    end else begin
      io_macOut = _27_19_inner_macOut;
    end
  end

  assign _zz__27_19_inner_macOut = ($signed(_zz__zz__27_19_inner_macOut) + $signed(_zz__zz__27_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_19_inner_activation <= 8'h00;
      _27_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_19_inner_activation <= io_addInput;
      end else begin
        _27_19_inner_macOut <= _zz__27_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_882 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_18_inner_macOut;
  wire       [15:0]   _zz__zz__27_18_inner_macOut_1;
  wire       [15:0]   _zz__27_18_inner_macOut_1;
  wire       [15:0]   _zz__27_18_inner_macOut_2;
  reg        [7:0]    _27_18_inner_activation;
  reg        [7:0]    _27_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_18_inner_macOut;

  assign _zz__zz__27_18_inner_macOut = ($signed(io_mulInput) * $signed(_27_18_inner_activation));
  assign _zz__zz__27_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_18_inner_macOut)) ? 16'h007f : _zz__27_18_inner_macOut_2);
  assign _zz__27_18_inner_macOut_2 = (($signed(_zz__27_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_18_inner_activation;
    end else begin
      io_macOut = _27_18_inner_macOut;
    end
  end

  assign _zz__27_18_inner_macOut = ($signed(_zz__zz__27_18_inner_macOut) + $signed(_zz__zz__27_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_18_inner_activation <= 8'h00;
      _27_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_18_inner_activation <= io_addInput;
      end else begin
        _27_18_inner_macOut <= _zz__27_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_881 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_17_inner_macOut;
  wire       [15:0]   _zz__zz__27_17_inner_macOut_1;
  wire       [15:0]   _zz__27_17_inner_macOut_1;
  wire       [15:0]   _zz__27_17_inner_macOut_2;
  reg        [7:0]    _27_17_inner_activation;
  reg        [7:0]    _27_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_17_inner_macOut;

  assign _zz__zz__27_17_inner_macOut = ($signed(io_mulInput) * $signed(_27_17_inner_activation));
  assign _zz__zz__27_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_17_inner_macOut)) ? 16'h007f : _zz__27_17_inner_macOut_2);
  assign _zz__27_17_inner_macOut_2 = (($signed(_zz__27_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_17_inner_activation;
    end else begin
      io_macOut = _27_17_inner_macOut;
    end
  end

  assign _zz__27_17_inner_macOut = ($signed(_zz__zz__27_17_inner_macOut) + $signed(_zz__zz__27_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_17_inner_activation <= 8'h00;
      _27_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_17_inner_activation <= io_addInput;
      end else begin
        _27_17_inner_macOut <= _zz__27_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_880 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_16_inner_macOut;
  wire       [15:0]   _zz__zz__27_16_inner_macOut_1;
  wire       [15:0]   _zz__27_16_inner_macOut_1;
  wire       [15:0]   _zz__27_16_inner_macOut_2;
  reg        [7:0]    _27_16_inner_activation;
  reg        [7:0]    _27_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_16_inner_macOut;

  assign _zz__zz__27_16_inner_macOut = ($signed(io_mulInput) * $signed(_27_16_inner_activation));
  assign _zz__zz__27_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_16_inner_macOut)) ? 16'h007f : _zz__27_16_inner_macOut_2);
  assign _zz__27_16_inner_macOut_2 = (($signed(_zz__27_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_16_inner_activation;
    end else begin
      io_macOut = _27_16_inner_macOut;
    end
  end

  assign _zz__27_16_inner_macOut = ($signed(_zz__zz__27_16_inner_macOut) + $signed(_zz__zz__27_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_16_inner_activation <= 8'h00;
      _27_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_16_inner_activation <= io_addInput;
      end else begin
        _27_16_inner_macOut <= _zz__27_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_879 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_15_inner_macOut;
  wire       [15:0]   _zz__zz__27_15_inner_macOut_1;
  wire       [15:0]   _zz__27_15_inner_macOut_1;
  wire       [15:0]   _zz__27_15_inner_macOut_2;
  reg        [7:0]    _27_15_inner_activation;
  reg        [7:0]    _27_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_15_inner_macOut;

  assign _zz__zz__27_15_inner_macOut = ($signed(io_mulInput) * $signed(_27_15_inner_activation));
  assign _zz__zz__27_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_15_inner_macOut)) ? 16'h007f : _zz__27_15_inner_macOut_2);
  assign _zz__27_15_inner_macOut_2 = (($signed(_zz__27_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_15_inner_activation;
    end else begin
      io_macOut = _27_15_inner_macOut;
    end
  end

  assign _zz__27_15_inner_macOut = ($signed(_zz__zz__27_15_inner_macOut) + $signed(_zz__zz__27_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_15_inner_activation <= 8'h00;
      _27_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_15_inner_activation <= io_addInput;
      end else begin
        _27_15_inner_macOut <= _zz__27_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_878 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_14_inner_macOut;
  wire       [15:0]   _zz__zz__27_14_inner_macOut_1;
  wire       [15:0]   _zz__27_14_inner_macOut_1;
  wire       [15:0]   _zz__27_14_inner_macOut_2;
  reg        [7:0]    _27_14_inner_activation;
  reg        [7:0]    _27_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_14_inner_macOut;

  assign _zz__zz__27_14_inner_macOut = ($signed(io_mulInput) * $signed(_27_14_inner_activation));
  assign _zz__zz__27_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_14_inner_macOut)) ? 16'h007f : _zz__27_14_inner_macOut_2);
  assign _zz__27_14_inner_macOut_2 = (($signed(_zz__27_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_14_inner_activation;
    end else begin
      io_macOut = _27_14_inner_macOut;
    end
  end

  assign _zz__27_14_inner_macOut = ($signed(_zz__zz__27_14_inner_macOut) + $signed(_zz__zz__27_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_14_inner_activation <= 8'h00;
      _27_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_14_inner_activation <= io_addInput;
      end else begin
        _27_14_inner_macOut <= _zz__27_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_877 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_13_inner_macOut;
  wire       [15:0]   _zz__zz__27_13_inner_macOut_1;
  wire       [15:0]   _zz__27_13_inner_macOut_1;
  wire       [15:0]   _zz__27_13_inner_macOut_2;
  reg        [7:0]    _27_13_inner_activation;
  reg        [7:0]    _27_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_13_inner_macOut;

  assign _zz__zz__27_13_inner_macOut = ($signed(io_mulInput) * $signed(_27_13_inner_activation));
  assign _zz__zz__27_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_13_inner_macOut)) ? 16'h007f : _zz__27_13_inner_macOut_2);
  assign _zz__27_13_inner_macOut_2 = (($signed(_zz__27_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_13_inner_activation;
    end else begin
      io_macOut = _27_13_inner_macOut;
    end
  end

  assign _zz__27_13_inner_macOut = ($signed(_zz__zz__27_13_inner_macOut) + $signed(_zz__zz__27_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_13_inner_activation <= 8'h00;
      _27_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_13_inner_activation <= io_addInput;
      end else begin
        _27_13_inner_macOut <= _zz__27_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_876 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_12_inner_macOut;
  wire       [15:0]   _zz__zz__27_12_inner_macOut_1;
  wire       [15:0]   _zz__27_12_inner_macOut_1;
  wire       [15:0]   _zz__27_12_inner_macOut_2;
  reg        [7:0]    _27_12_inner_activation;
  reg        [7:0]    _27_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_12_inner_macOut;

  assign _zz__zz__27_12_inner_macOut = ($signed(io_mulInput) * $signed(_27_12_inner_activation));
  assign _zz__zz__27_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_12_inner_macOut)) ? 16'h007f : _zz__27_12_inner_macOut_2);
  assign _zz__27_12_inner_macOut_2 = (($signed(_zz__27_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_12_inner_activation;
    end else begin
      io_macOut = _27_12_inner_macOut;
    end
  end

  assign _zz__27_12_inner_macOut = ($signed(_zz__zz__27_12_inner_macOut) + $signed(_zz__zz__27_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_12_inner_activation <= 8'h00;
      _27_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_12_inner_activation <= io_addInput;
      end else begin
        _27_12_inner_macOut <= _zz__27_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_875 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_11_inner_macOut;
  wire       [15:0]   _zz__zz__27_11_inner_macOut_1;
  wire       [15:0]   _zz__27_11_inner_macOut_1;
  wire       [15:0]   _zz__27_11_inner_macOut_2;
  reg        [7:0]    _27_11_inner_activation;
  reg        [7:0]    _27_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_11_inner_macOut;

  assign _zz__zz__27_11_inner_macOut = ($signed(io_mulInput) * $signed(_27_11_inner_activation));
  assign _zz__zz__27_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_11_inner_macOut)) ? 16'h007f : _zz__27_11_inner_macOut_2);
  assign _zz__27_11_inner_macOut_2 = (($signed(_zz__27_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_11_inner_activation;
    end else begin
      io_macOut = _27_11_inner_macOut;
    end
  end

  assign _zz__27_11_inner_macOut = ($signed(_zz__zz__27_11_inner_macOut) + $signed(_zz__zz__27_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_11_inner_activation <= 8'h00;
      _27_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_11_inner_activation <= io_addInput;
      end else begin
        _27_11_inner_macOut <= _zz__27_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_874 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_10_inner_macOut;
  wire       [15:0]   _zz__zz__27_10_inner_macOut_1;
  wire       [15:0]   _zz__27_10_inner_macOut_1;
  wire       [15:0]   _zz__27_10_inner_macOut_2;
  reg        [7:0]    _27_10_inner_activation;
  reg        [7:0]    _27_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_10_inner_macOut;

  assign _zz__zz__27_10_inner_macOut = ($signed(io_mulInput) * $signed(_27_10_inner_activation));
  assign _zz__zz__27_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_10_inner_macOut)) ? 16'h007f : _zz__27_10_inner_macOut_2);
  assign _zz__27_10_inner_macOut_2 = (($signed(_zz__27_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_10_inner_activation;
    end else begin
      io_macOut = _27_10_inner_macOut;
    end
  end

  assign _zz__27_10_inner_macOut = ($signed(_zz__zz__27_10_inner_macOut) + $signed(_zz__zz__27_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_10_inner_activation <= 8'h00;
      _27_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_10_inner_activation <= io_addInput;
      end else begin
        _27_10_inner_macOut <= _zz__27_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_873 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_9_inner_macOut;
  wire       [15:0]   _zz__zz__27_9_inner_macOut_1;
  wire       [15:0]   _zz__27_9_inner_macOut_1;
  wire       [15:0]   _zz__27_9_inner_macOut_2;
  reg        [7:0]    _27_9_inner_activation;
  reg        [7:0]    _27_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_9_inner_macOut;

  assign _zz__zz__27_9_inner_macOut = ($signed(io_mulInput) * $signed(_27_9_inner_activation));
  assign _zz__zz__27_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_9_inner_macOut)) ? 16'h007f : _zz__27_9_inner_macOut_2);
  assign _zz__27_9_inner_macOut_2 = (($signed(_zz__27_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_9_inner_activation;
    end else begin
      io_macOut = _27_9_inner_macOut;
    end
  end

  assign _zz__27_9_inner_macOut = ($signed(_zz__zz__27_9_inner_macOut) + $signed(_zz__zz__27_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_9_inner_activation <= 8'h00;
      _27_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_9_inner_activation <= io_addInput;
      end else begin
        _27_9_inner_macOut <= _zz__27_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_872 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_8_inner_macOut;
  wire       [15:0]   _zz__zz__27_8_inner_macOut_1;
  wire       [15:0]   _zz__27_8_inner_macOut_1;
  wire       [15:0]   _zz__27_8_inner_macOut_2;
  reg        [7:0]    _27_8_inner_activation;
  reg        [7:0]    _27_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_8_inner_macOut;

  assign _zz__zz__27_8_inner_macOut = ($signed(io_mulInput) * $signed(_27_8_inner_activation));
  assign _zz__zz__27_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_8_inner_macOut)) ? 16'h007f : _zz__27_8_inner_macOut_2);
  assign _zz__27_8_inner_macOut_2 = (($signed(_zz__27_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_8_inner_activation;
    end else begin
      io_macOut = _27_8_inner_macOut;
    end
  end

  assign _zz__27_8_inner_macOut = ($signed(_zz__zz__27_8_inner_macOut) + $signed(_zz__zz__27_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_8_inner_activation <= 8'h00;
      _27_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_8_inner_activation <= io_addInput;
      end else begin
        _27_8_inner_macOut <= _zz__27_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_871 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_7_inner_macOut;
  wire       [15:0]   _zz__zz__27_7_inner_macOut_1;
  wire       [15:0]   _zz__27_7_inner_macOut_1;
  wire       [15:0]   _zz__27_7_inner_macOut_2;
  reg        [7:0]    _27_7_inner_activation;
  reg        [7:0]    _27_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_7_inner_macOut;

  assign _zz__zz__27_7_inner_macOut = ($signed(io_mulInput) * $signed(_27_7_inner_activation));
  assign _zz__zz__27_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_7_inner_macOut)) ? 16'h007f : _zz__27_7_inner_macOut_2);
  assign _zz__27_7_inner_macOut_2 = (($signed(_zz__27_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_7_inner_activation;
    end else begin
      io_macOut = _27_7_inner_macOut;
    end
  end

  assign _zz__27_7_inner_macOut = ($signed(_zz__zz__27_7_inner_macOut) + $signed(_zz__zz__27_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_7_inner_activation <= 8'h00;
      _27_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_7_inner_activation <= io_addInput;
      end else begin
        _27_7_inner_macOut <= _zz__27_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_870 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_6_inner_macOut;
  wire       [15:0]   _zz__zz__27_6_inner_macOut_1;
  wire       [15:0]   _zz__27_6_inner_macOut_1;
  wire       [15:0]   _zz__27_6_inner_macOut_2;
  reg        [7:0]    _27_6_inner_activation;
  reg        [7:0]    _27_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_6_inner_macOut;

  assign _zz__zz__27_6_inner_macOut = ($signed(io_mulInput) * $signed(_27_6_inner_activation));
  assign _zz__zz__27_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_6_inner_macOut)) ? 16'h007f : _zz__27_6_inner_macOut_2);
  assign _zz__27_6_inner_macOut_2 = (($signed(_zz__27_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_6_inner_activation;
    end else begin
      io_macOut = _27_6_inner_macOut;
    end
  end

  assign _zz__27_6_inner_macOut = ($signed(_zz__zz__27_6_inner_macOut) + $signed(_zz__zz__27_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_6_inner_activation <= 8'h00;
      _27_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_6_inner_activation <= io_addInput;
      end else begin
        _27_6_inner_macOut <= _zz__27_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_869 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_5_inner_macOut;
  wire       [15:0]   _zz__zz__27_5_inner_macOut_1;
  wire       [15:0]   _zz__27_5_inner_macOut_1;
  wire       [15:0]   _zz__27_5_inner_macOut_2;
  reg        [7:0]    _27_5_inner_activation;
  reg        [7:0]    _27_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_5_inner_macOut;

  assign _zz__zz__27_5_inner_macOut = ($signed(io_mulInput) * $signed(_27_5_inner_activation));
  assign _zz__zz__27_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_5_inner_macOut)) ? 16'h007f : _zz__27_5_inner_macOut_2);
  assign _zz__27_5_inner_macOut_2 = (($signed(_zz__27_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_5_inner_activation;
    end else begin
      io_macOut = _27_5_inner_macOut;
    end
  end

  assign _zz__27_5_inner_macOut = ($signed(_zz__zz__27_5_inner_macOut) + $signed(_zz__zz__27_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_5_inner_activation <= 8'h00;
      _27_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_5_inner_activation <= io_addInput;
      end else begin
        _27_5_inner_macOut <= _zz__27_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_868 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_4_inner_macOut;
  wire       [15:0]   _zz__zz__27_4_inner_macOut_1;
  wire       [15:0]   _zz__27_4_inner_macOut_1;
  wire       [15:0]   _zz__27_4_inner_macOut_2;
  reg        [7:0]    _27_4_inner_activation;
  reg        [7:0]    _27_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_4_inner_macOut;

  assign _zz__zz__27_4_inner_macOut = ($signed(io_mulInput) * $signed(_27_4_inner_activation));
  assign _zz__zz__27_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_4_inner_macOut)) ? 16'h007f : _zz__27_4_inner_macOut_2);
  assign _zz__27_4_inner_macOut_2 = (($signed(_zz__27_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_4_inner_activation;
    end else begin
      io_macOut = _27_4_inner_macOut;
    end
  end

  assign _zz__27_4_inner_macOut = ($signed(_zz__zz__27_4_inner_macOut) + $signed(_zz__zz__27_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_4_inner_activation <= 8'h00;
      _27_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_4_inner_activation <= io_addInput;
      end else begin
        _27_4_inner_macOut <= _zz__27_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_867 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_3_inner_macOut;
  wire       [15:0]   _zz__zz__27_3_inner_macOut_1;
  wire       [15:0]   _zz__27_3_inner_macOut_1;
  wire       [15:0]   _zz__27_3_inner_macOut_2;
  reg        [7:0]    _27_3_inner_activation;
  reg        [7:0]    _27_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_3_inner_macOut;

  assign _zz__zz__27_3_inner_macOut = ($signed(io_mulInput) * $signed(_27_3_inner_activation));
  assign _zz__zz__27_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_3_inner_macOut)) ? 16'h007f : _zz__27_3_inner_macOut_2);
  assign _zz__27_3_inner_macOut_2 = (($signed(_zz__27_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_3_inner_activation;
    end else begin
      io_macOut = _27_3_inner_macOut;
    end
  end

  assign _zz__27_3_inner_macOut = ($signed(_zz__zz__27_3_inner_macOut) + $signed(_zz__zz__27_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_3_inner_activation <= 8'h00;
      _27_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_3_inner_activation <= io_addInput;
      end else begin
        _27_3_inner_macOut <= _zz__27_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_866 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_2_inner_macOut;
  wire       [15:0]   _zz__zz__27_2_inner_macOut_1;
  wire       [15:0]   _zz__27_2_inner_macOut_1;
  wire       [15:0]   _zz__27_2_inner_macOut_2;
  reg        [7:0]    _27_2_inner_activation;
  reg        [7:0]    _27_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_2_inner_macOut;

  assign _zz__zz__27_2_inner_macOut = ($signed(io_mulInput) * $signed(_27_2_inner_activation));
  assign _zz__zz__27_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_2_inner_macOut)) ? 16'h007f : _zz__27_2_inner_macOut_2);
  assign _zz__27_2_inner_macOut_2 = (($signed(_zz__27_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_2_inner_activation;
    end else begin
      io_macOut = _27_2_inner_macOut;
    end
  end

  assign _zz__27_2_inner_macOut = ($signed(_zz__zz__27_2_inner_macOut) + $signed(_zz__zz__27_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_2_inner_activation <= 8'h00;
      _27_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_2_inner_activation <= io_addInput;
      end else begin
        _27_2_inner_macOut <= _zz__27_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_865 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_1_inner_macOut;
  wire       [15:0]   _zz__zz__27_1_inner_macOut_1;
  wire       [15:0]   _zz__27_1_inner_macOut_1;
  wire       [15:0]   _zz__27_1_inner_macOut_2;
  reg        [7:0]    _27_1_inner_activation;
  reg        [7:0]    _27_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_1_inner_macOut;

  assign _zz__zz__27_1_inner_macOut = ($signed(io_mulInput) * $signed(_27_1_inner_activation));
  assign _zz__zz__27_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_1_inner_macOut)) ? 16'h007f : _zz__27_1_inner_macOut_2);
  assign _zz__27_1_inner_macOut_2 = (($signed(_zz__27_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_1_inner_activation;
    end else begin
      io_macOut = _27_1_inner_macOut;
    end
  end

  assign _zz__27_1_inner_macOut = ($signed(_zz__zz__27_1_inner_macOut) + $signed(_zz__zz__27_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_1_inner_activation <= 8'h00;
      _27_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_1_inner_activation <= io_addInput;
      end else begin
        _27_1_inner_macOut <= _zz__27_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_864 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__27_0_inner_macOut;
  wire       [15:0]   _zz__zz__27_0_inner_macOut_1;
  wire       [15:0]   _zz__27_0_inner_macOut_1;
  wire       [15:0]   _zz__27_0_inner_macOut_2;
  reg        [7:0]    _27_0_inner_activation;
  reg        [7:0]    _27_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__27_0_inner_macOut;

  assign _zz__zz__27_0_inner_macOut = ($signed(io_mulInput) * $signed(_27_0_inner_activation));
  assign _zz__zz__27_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__27_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__27_0_inner_macOut)) ? 16'h007f : _zz__27_0_inner_macOut_2);
  assign _zz__27_0_inner_macOut_2 = (($signed(_zz__27_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__27_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _27_0_inner_activation;
    end else begin
      io_macOut = _27_0_inner_macOut;
    end
  end

  assign _zz__27_0_inner_macOut = ($signed(_zz__zz__27_0_inner_macOut) + $signed(_zz__zz__27_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _27_0_inner_activation <= 8'h00;
      _27_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _27_0_inner_activation <= io_addInput;
      end else begin
        _27_0_inner_macOut <= _zz__27_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_863 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_31_inner_macOut;
  wire       [15:0]   _zz__zz__26_31_inner_macOut_1;
  wire       [15:0]   _zz__26_31_inner_macOut_1;
  wire       [15:0]   _zz__26_31_inner_macOut_2;
  reg        [7:0]    _26_31_inner_activation;
  reg        [7:0]    _26_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_31_inner_macOut;

  assign _zz__zz__26_31_inner_macOut = ($signed(io_mulInput) * $signed(_26_31_inner_activation));
  assign _zz__zz__26_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_31_inner_macOut)) ? 16'h007f : _zz__26_31_inner_macOut_2);
  assign _zz__26_31_inner_macOut_2 = (($signed(_zz__26_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_31_inner_activation;
    end else begin
      io_macOut = _26_31_inner_macOut;
    end
  end

  assign _zz__26_31_inner_macOut = ($signed(_zz__zz__26_31_inner_macOut) + $signed(_zz__zz__26_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_31_inner_activation <= 8'h00;
      _26_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_31_inner_activation <= io_addInput;
      end else begin
        _26_31_inner_macOut <= _zz__26_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_862 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_30_inner_macOut;
  wire       [15:0]   _zz__zz__26_30_inner_macOut_1;
  wire       [15:0]   _zz__26_30_inner_macOut_1;
  wire       [15:0]   _zz__26_30_inner_macOut_2;
  reg        [7:0]    _26_30_inner_activation;
  reg        [7:0]    _26_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_30_inner_macOut;

  assign _zz__zz__26_30_inner_macOut = ($signed(io_mulInput) * $signed(_26_30_inner_activation));
  assign _zz__zz__26_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_30_inner_macOut)) ? 16'h007f : _zz__26_30_inner_macOut_2);
  assign _zz__26_30_inner_macOut_2 = (($signed(_zz__26_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_30_inner_activation;
    end else begin
      io_macOut = _26_30_inner_macOut;
    end
  end

  assign _zz__26_30_inner_macOut = ($signed(_zz__zz__26_30_inner_macOut) + $signed(_zz__zz__26_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_30_inner_activation <= 8'h00;
      _26_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_30_inner_activation <= io_addInput;
      end else begin
        _26_30_inner_macOut <= _zz__26_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_861 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_29_inner_macOut;
  wire       [15:0]   _zz__zz__26_29_inner_macOut_1;
  wire       [15:0]   _zz__26_29_inner_macOut_1;
  wire       [15:0]   _zz__26_29_inner_macOut_2;
  reg        [7:0]    _26_29_inner_activation;
  reg        [7:0]    _26_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_29_inner_macOut;

  assign _zz__zz__26_29_inner_macOut = ($signed(io_mulInput) * $signed(_26_29_inner_activation));
  assign _zz__zz__26_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_29_inner_macOut)) ? 16'h007f : _zz__26_29_inner_macOut_2);
  assign _zz__26_29_inner_macOut_2 = (($signed(_zz__26_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_29_inner_activation;
    end else begin
      io_macOut = _26_29_inner_macOut;
    end
  end

  assign _zz__26_29_inner_macOut = ($signed(_zz__zz__26_29_inner_macOut) + $signed(_zz__zz__26_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_29_inner_activation <= 8'h00;
      _26_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_29_inner_activation <= io_addInput;
      end else begin
        _26_29_inner_macOut <= _zz__26_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_860 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_28_inner_macOut;
  wire       [15:0]   _zz__zz__26_28_inner_macOut_1;
  wire       [15:0]   _zz__26_28_inner_macOut_1;
  wire       [15:0]   _zz__26_28_inner_macOut_2;
  reg        [7:0]    _26_28_inner_activation;
  reg        [7:0]    _26_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_28_inner_macOut;

  assign _zz__zz__26_28_inner_macOut = ($signed(io_mulInput) * $signed(_26_28_inner_activation));
  assign _zz__zz__26_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_28_inner_macOut)) ? 16'h007f : _zz__26_28_inner_macOut_2);
  assign _zz__26_28_inner_macOut_2 = (($signed(_zz__26_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_28_inner_activation;
    end else begin
      io_macOut = _26_28_inner_macOut;
    end
  end

  assign _zz__26_28_inner_macOut = ($signed(_zz__zz__26_28_inner_macOut) + $signed(_zz__zz__26_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_28_inner_activation <= 8'h00;
      _26_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_28_inner_activation <= io_addInput;
      end else begin
        _26_28_inner_macOut <= _zz__26_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_859 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_27_inner_macOut;
  wire       [15:0]   _zz__zz__26_27_inner_macOut_1;
  wire       [15:0]   _zz__26_27_inner_macOut_1;
  wire       [15:0]   _zz__26_27_inner_macOut_2;
  reg        [7:0]    _26_27_inner_activation;
  reg        [7:0]    _26_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_27_inner_macOut;

  assign _zz__zz__26_27_inner_macOut = ($signed(io_mulInput) * $signed(_26_27_inner_activation));
  assign _zz__zz__26_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_27_inner_macOut)) ? 16'h007f : _zz__26_27_inner_macOut_2);
  assign _zz__26_27_inner_macOut_2 = (($signed(_zz__26_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_27_inner_activation;
    end else begin
      io_macOut = _26_27_inner_macOut;
    end
  end

  assign _zz__26_27_inner_macOut = ($signed(_zz__zz__26_27_inner_macOut) + $signed(_zz__zz__26_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_27_inner_activation <= 8'h00;
      _26_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_27_inner_activation <= io_addInput;
      end else begin
        _26_27_inner_macOut <= _zz__26_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_858 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_26_inner_macOut;
  wire       [15:0]   _zz__zz__26_26_inner_macOut_1;
  wire       [15:0]   _zz__26_26_inner_macOut_1;
  wire       [15:0]   _zz__26_26_inner_macOut_2;
  reg        [7:0]    _26_26_inner_activation;
  reg        [7:0]    _26_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_26_inner_macOut;

  assign _zz__zz__26_26_inner_macOut = ($signed(io_mulInput) * $signed(_26_26_inner_activation));
  assign _zz__zz__26_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_26_inner_macOut)) ? 16'h007f : _zz__26_26_inner_macOut_2);
  assign _zz__26_26_inner_macOut_2 = (($signed(_zz__26_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_26_inner_activation;
    end else begin
      io_macOut = _26_26_inner_macOut;
    end
  end

  assign _zz__26_26_inner_macOut = ($signed(_zz__zz__26_26_inner_macOut) + $signed(_zz__zz__26_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_26_inner_activation <= 8'h00;
      _26_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_26_inner_activation <= io_addInput;
      end else begin
        _26_26_inner_macOut <= _zz__26_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_857 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_25_inner_macOut;
  wire       [15:0]   _zz__zz__26_25_inner_macOut_1;
  wire       [15:0]   _zz__26_25_inner_macOut_1;
  wire       [15:0]   _zz__26_25_inner_macOut_2;
  reg        [7:0]    _26_25_inner_activation;
  reg        [7:0]    _26_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_25_inner_macOut;

  assign _zz__zz__26_25_inner_macOut = ($signed(io_mulInput) * $signed(_26_25_inner_activation));
  assign _zz__zz__26_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_25_inner_macOut)) ? 16'h007f : _zz__26_25_inner_macOut_2);
  assign _zz__26_25_inner_macOut_2 = (($signed(_zz__26_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_25_inner_activation;
    end else begin
      io_macOut = _26_25_inner_macOut;
    end
  end

  assign _zz__26_25_inner_macOut = ($signed(_zz__zz__26_25_inner_macOut) + $signed(_zz__zz__26_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_25_inner_activation <= 8'h00;
      _26_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_25_inner_activation <= io_addInput;
      end else begin
        _26_25_inner_macOut <= _zz__26_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_856 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_24_inner_macOut;
  wire       [15:0]   _zz__zz__26_24_inner_macOut_1;
  wire       [15:0]   _zz__26_24_inner_macOut_1;
  wire       [15:0]   _zz__26_24_inner_macOut_2;
  reg        [7:0]    _26_24_inner_activation;
  reg        [7:0]    _26_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_24_inner_macOut;

  assign _zz__zz__26_24_inner_macOut = ($signed(io_mulInput) * $signed(_26_24_inner_activation));
  assign _zz__zz__26_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_24_inner_macOut)) ? 16'h007f : _zz__26_24_inner_macOut_2);
  assign _zz__26_24_inner_macOut_2 = (($signed(_zz__26_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_24_inner_activation;
    end else begin
      io_macOut = _26_24_inner_macOut;
    end
  end

  assign _zz__26_24_inner_macOut = ($signed(_zz__zz__26_24_inner_macOut) + $signed(_zz__zz__26_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_24_inner_activation <= 8'h00;
      _26_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_24_inner_activation <= io_addInput;
      end else begin
        _26_24_inner_macOut <= _zz__26_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_855 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_23_inner_macOut;
  wire       [15:0]   _zz__zz__26_23_inner_macOut_1;
  wire       [15:0]   _zz__26_23_inner_macOut_1;
  wire       [15:0]   _zz__26_23_inner_macOut_2;
  reg        [7:0]    _26_23_inner_activation;
  reg        [7:0]    _26_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_23_inner_macOut;

  assign _zz__zz__26_23_inner_macOut = ($signed(io_mulInput) * $signed(_26_23_inner_activation));
  assign _zz__zz__26_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_23_inner_macOut)) ? 16'h007f : _zz__26_23_inner_macOut_2);
  assign _zz__26_23_inner_macOut_2 = (($signed(_zz__26_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_23_inner_activation;
    end else begin
      io_macOut = _26_23_inner_macOut;
    end
  end

  assign _zz__26_23_inner_macOut = ($signed(_zz__zz__26_23_inner_macOut) + $signed(_zz__zz__26_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_23_inner_activation <= 8'h00;
      _26_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_23_inner_activation <= io_addInput;
      end else begin
        _26_23_inner_macOut <= _zz__26_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_854 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_22_inner_macOut;
  wire       [15:0]   _zz__zz__26_22_inner_macOut_1;
  wire       [15:0]   _zz__26_22_inner_macOut_1;
  wire       [15:0]   _zz__26_22_inner_macOut_2;
  reg        [7:0]    _26_22_inner_activation;
  reg        [7:0]    _26_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_22_inner_macOut;

  assign _zz__zz__26_22_inner_macOut = ($signed(io_mulInput) * $signed(_26_22_inner_activation));
  assign _zz__zz__26_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_22_inner_macOut)) ? 16'h007f : _zz__26_22_inner_macOut_2);
  assign _zz__26_22_inner_macOut_2 = (($signed(_zz__26_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_22_inner_activation;
    end else begin
      io_macOut = _26_22_inner_macOut;
    end
  end

  assign _zz__26_22_inner_macOut = ($signed(_zz__zz__26_22_inner_macOut) + $signed(_zz__zz__26_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_22_inner_activation <= 8'h00;
      _26_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_22_inner_activation <= io_addInput;
      end else begin
        _26_22_inner_macOut <= _zz__26_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_853 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_21_inner_macOut;
  wire       [15:0]   _zz__zz__26_21_inner_macOut_1;
  wire       [15:0]   _zz__26_21_inner_macOut_1;
  wire       [15:0]   _zz__26_21_inner_macOut_2;
  reg        [7:0]    _26_21_inner_activation;
  reg        [7:0]    _26_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_21_inner_macOut;

  assign _zz__zz__26_21_inner_macOut = ($signed(io_mulInput) * $signed(_26_21_inner_activation));
  assign _zz__zz__26_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_21_inner_macOut)) ? 16'h007f : _zz__26_21_inner_macOut_2);
  assign _zz__26_21_inner_macOut_2 = (($signed(_zz__26_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_21_inner_activation;
    end else begin
      io_macOut = _26_21_inner_macOut;
    end
  end

  assign _zz__26_21_inner_macOut = ($signed(_zz__zz__26_21_inner_macOut) + $signed(_zz__zz__26_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_21_inner_activation <= 8'h00;
      _26_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_21_inner_activation <= io_addInput;
      end else begin
        _26_21_inner_macOut <= _zz__26_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_852 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_20_inner_macOut;
  wire       [15:0]   _zz__zz__26_20_inner_macOut_1;
  wire       [15:0]   _zz__26_20_inner_macOut_1;
  wire       [15:0]   _zz__26_20_inner_macOut_2;
  reg        [7:0]    _26_20_inner_activation;
  reg        [7:0]    _26_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_20_inner_macOut;

  assign _zz__zz__26_20_inner_macOut = ($signed(io_mulInput) * $signed(_26_20_inner_activation));
  assign _zz__zz__26_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_20_inner_macOut)) ? 16'h007f : _zz__26_20_inner_macOut_2);
  assign _zz__26_20_inner_macOut_2 = (($signed(_zz__26_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_20_inner_activation;
    end else begin
      io_macOut = _26_20_inner_macOut;
    end
  end

  assign _zz__26_20_inner_macOut = ($signed(_zz__zz__26_20_inner_macOut) + $signed(_zz__zz__26_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_20_inner_activation <= 8'h00;
      _26_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_20_inner_activation <= io_addInput;
      end else begin
        _26_20_inner_macOut <= _zz__26_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_851 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_19_inner_macOut;
  wire       [15:0]   _zz__zz__26_19_inner_macOut_1;
  wire       [15:0]   _zz__26_19_inner_macOut_1;
  wire       [15:0]   _zz__26_19_inner_macOut_2;
  reg        [7:0]    _26_19_inner_activation;
  reg        [7:0]    _26_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_19_inner_macOut;

  assign _zz__zz__26_19_inner_macOut = ($signed(io_mulInput) * $signed(_26_19_inner_activation));
  assign _zz__zz__26_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_19_inner_macOut)) ? 16'h007f : _zz__26_19_inner_macOut_2);
  assign _zz__26_19_inner_macOut_2 = (($signed(_zz__26_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_19_inner_activation;
    end else begin
      io_macOut = _26_19_inner_macOut;
    end
  end

  assign _zz__26_19_inner_macOut = ($signed(_zz__zz__26_19_inner_macOut) + $signed(_zz__zz__26_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_19_inner_activation <= 8'h00;
      _26_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_19_inner_activation <= io_addInput;
      end else begin
        _26_19_inner_macOut <= _zz__26_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_850 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_18_inner_macOut;
  wire       [15:0]   _zz__zz__26_18_inner_macOut_1;
  wire       [15:0]   _zz__26_18_inner_macOut_1;
  wire       [15:0]   _zz__26_18_inner_macOut_2;
  reg        [7:0]    _26_18_inner_activation;
  reg        [7:0]    _26_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_18_inner_macOut;

  assign _zz__zz__26_18_inner_macOut = ($signed(io_mulInput) * $signed(_26_18_inner_activation));
  assign _zz__zz__26_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_18_inner_macOut)) ? 16'h007f : _zz__26_18_inner_macOut_2);
  assign _zz__26_18_inner_macOut_2 = (($signed(_zz__26_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_18_inner_activation;
    end else begin
      io_macOut = _26_18_inner_macOut;
    end
  end

  assign _zz__26_18_inner_macOut = ($signed(_zz__zz__26_18_inner_macOut) + $signed(_zz__zz__26_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_18_inner_activation <= 8'h00;
      _26_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_18_inner_activation <= io_addInput;
      end else begin
        _26_18_inner_macOut <= _zz__26_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_849 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_17_inner_macOut;
  wire       [15:0]   _zz__zz__26_17_inner_macOut_1;
  wire       [15:0]   _zz__26_17_inner_macOut_1;
  wire       [15:0]   _zz__26_17_inner_macOut_2;
  reg        [7:0]    _26_17_inner_activation;
  reg        [7:0]    _26_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_17_inner_macOut;

  assign _zz__zz__26_17_inner_macOut = ($signed(io_mulInput) * $signed(_26_17_inner_activation));
  assign _zz__zz__26_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_17_inner_macOut)) ? 16'h007f : _zz__26_17_inner_macOut_2);
  assign _zz__26_17_inner_macOut_2 = (($signed(_zz__26_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_17_inner_activation;
    end else begin
      io_macOut = _26_17_inner_macOut;
    end
  end

  assign _zz__26_17_inner_macOut = ($signed(_zz__zz__26_17_inner_macOut) + $signed(_zz__zz__26_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_17_inner_activation <= 8'h00;
      _26_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_17_inner_activation <= io_addInput;
      end else begin
        _26_17_inner_macOut <= _zz__26_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_848 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_16_inner_macOut;
  wire       [15:0]   _zz__zz__26_16_inner_macOut_1;
  wire       [15:0]   _zz__26_16_inner_macOut_1;
  wire       [15:0]   _zz__26_16_inner_macOut_2;
  reg        [7:0]    _26_16_inner_activation;
  reg        [7:0]    _26_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_16_inner_macOut;

  assign _zz__zz__26_16_inner_macOut = ($signed(io_mulInput) * $signed(_26_16_inner_activation));
  assign _zz__zz__26_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_16_inner_macOut)) ? 16'h007f : _zz__26_16_inner_macOut_2);
  assign _zz__26_16_inner_macOut_2 = (($signed(_zz__26_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_16_inner_activation;
    end else begin
      io_macOut = _26_16_inner_macOut;
    end
  end

  assign _zz__26_16_inner_macOut = ($signed(_zz__zz__26_16_inner_macOut) + $signed(_zz__zz__26_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_16_inner_activation <= 8'h00;
      _26_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_16_inner_activation <= io_addInput;
      end else begin
        _26_16_inner_macOut <= _zz__26_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_847 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_15_inner_macOut;
  wire       [15:0]   _zz__zz__26_15_inner_macOut_1;
  wire       [15:0]   _zz__26_15_inner_macOut_1;
  wire       [15:0]   _zz__26_15_inner_macOut_2;
  reg        [7:0]    _26_15_inner_activation;
  reg        [7:0]    _26_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_15_inner_macOut;

  assign _zz__zz__26_15_inner_macOut = ($signed(io_mulInput) * $signed(_26_15_inner_activation));
  assign _zz__zz__26_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_15_inner_macOut)) ? 16'h007f : _zz__26_15_inner_macOut_2);
  assign _zz__26_15_inner_macOut_2 = (($signed(_zz__26_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_15_inner_activation;
    end else begin
      io_macOut = _26_15_inner_macOut;
    end
  end

  assign _zz__26_15_inner_macOut = ($signed(_zz__zz__26_15_inner_macOut) + $signed(_zz__zz__26_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_15_inner_activation <= 8'h00;
      _26_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_15_inner_activation <= io_addInput;
      end else begin
        _26_15_inner_macOut <= _zz__26_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_846 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_14_inner_macOut;
  wire       [15:0]   _zz__zz__26_14_inner_macOut_1;
  wire       [15:0]   _zz__26_14_inner_macOut_1;
  wire       [15:0]   _zz__26_14_inner_macOut_2;
  reg        [7:0]    _26_14_inner_activation;
  reg        [7:0]    _26_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_14_inner_macOut;

  assign _zz__zz__26_14_inner_macOut = ($signed(io_mulInput) * $signed(_26_14_inner_activation));
  assign _zz__zz__26_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_14_inner_macOut)) ? 16'h007f : _zz__26_14_inner_macOut_2);
  assign _zz__26_14_inner_macOut_2 = (($signed(_zz__26_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_14_inner_activation;
    end else begin
      io_macOut = _26_14_inner_macOut;
    end
  end

  assign _zz__26_14_inner_macOut = ($signed(_zz__zz__26_14_inner_macOut) + $signed(_zz__zz__26_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_14_inner_activation <= 8'h00;
      _26_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_14_inner_activation <= io_addInput;
      end else begin
        _26_14_inner_macOut <= _zz__26_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_845 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_13_inner_macOut;
  wire       [15:0]   _zz__zz__26_13_inner_macOut_1;
  wire       [15:0]   _zz__26_13_inner_macOut_1;
  wire       [15:0]   _zz__26_13_inner_macOut_2;
  reg        [7:0]    _26_13_inner_activation;
  reg        [7:0]    _26_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_13_inner_macOut;

  assign _zz__zz__26_13_inner_macOut = ($signed(io_mulInput) * $signed(_26_13_inner_activation));
  assign _zz__zz__26_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_13_inner_macOut)) ? 16'h007f : _zz__26_13_inner_macOut_2);
  assign _zz__26_13_inner_macOut_2 = (($signed(_zz__26_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_13_inner_activation;
    end else begin
      io_macOut = _26_13_inner_macOut;
    end
  end

  assign _zz__26_13_inner_macOut = ($signed(_zz__zz__26_13_inner_macOut) + $signed(_zz__zz__26_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_13_inner_activation <= 8'h00;
      _26_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_13_inner_activation <= io_addInput;
      end else begin
        _26_13_inner_macOut <= _zz__26_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_844 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_12_inner_macOut;
  wire       [15:0]   _zz__zz__26_12_inner_macOut_1;
  wire       [15:0]   _zz__26_12_inner_macOut_1;
  wire       [15:0]   _zz__26_12_inner_macOut_2;
  reg        [7:0]    _26_12_inner_activation;
  reg        [7:0]    _26_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_12_inner_macOut;

  assign _zz__zz__26_12_inner_macOut = ($signed(io_mulInput) * $signed(_26_12_inner_activation));
  assign _zz__zz__26_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_12_inner_macOut)) ? 16'h007f : _zz__26_12_inner_macOut_2);
  assign _zz__26_12_inner_macOut_2 = (($signed(_zz__26_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_12_inner_activation;
    end else begin
      io_macOut = _26_12_inner_macOut;
    end
  end

  assign _zz__26_12_inner_macOut = ($signed(_zz__zz__26_12_inner_macOut) + $signed(_zz__zz__26_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_12_inner_activation <= 8'h00;
      _26_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_12_inner_activation <= io_addInput;
      end else begin
        _26_12_inner_macOut <= _zz__26_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_843 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_11_inner_macOut;
  wire       [15:0]   _zz__zz__26_11_inner_macOut_1;
  wire       [15:0]   _zz__26_11_inner_macOut_1;
  wire       [15:0]   _zz__26_11_inner_macOut_2;
  reg        [7:0]    _26_11_inner_activation;
  reg        [7:0]    _26_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_11_inner_macOut;

  assign _zz__zz__26_11_inner_macOut = ($signed(io_mulInput) * $signed(_26_11_inner_activation));
  assign _zz__zz__26_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_11_inner_macOut)) ? 16'h007f : _zz__26_11_inner_macOut_2);
  assign _zz__26_11_inner_macOut_2 = (($signed(_zz__26_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_11_inner_activation;
    end else begin
      io_macOut = _26_11_inner_macOut;
    end
  end

  assign _zz__26_11_inner_macOut = ($signed(_zz__zz__26_11_inner_macOut) + $signed(_zz__zz__26_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_11_inner_activation <= 8'h00;
      _26_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_11_inner_activation <= io_addInput;
      end else begin
        _26_11_inner_macOut <= _zz__26_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_842 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_10_inner_macOut;
  wire       [15:0]   _zz__zz__26_10_inner_macOut_1;
  wire       [15:0]   _zz__26_10_inner_macOut_1;
  wire       [15:0]   _zz__26_10_inner_macOut_2;
  reg        [7:0]    _26_10_inner_activation;
  reg        [7:0]    _26_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_10_inner_macOut;

  assign _zz__zz__26_10_inner_macOut = ($signed(io_mulInput) * $signed(_26_10_inner_activation));
  assign _zz__zz__26_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_10_inner_macOut)) ? 16'h007f : _zz__26_10_inner_macOut_2);
  assign _zz__26_10_inner_macOut_2 = (($signed(_zz__26_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_10_inner_activation;
    end else begin
      io_macOut = _26_10_inner_macOut;
    end
  end

  assign _zz__26_10_inner_macOut = ($signed(_zz__zz__26_10_inner_macOut) + $signed(_zz__zz__26_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_10_inner_activation <= 8'h00;
      _26_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_10_inner_activation <= io_addInput;
      end else begin
        _26_10_inner_macOut <= _zz__26_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_841 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_9_inner_macOut;
  wire       [15:0]   _zz__zz__26_9_inner_macOut_1;
  wire       [15:0]   _zz__26_9_inner_macOut_1;
  wire       [15:0]   _zz__26_9_inner_macOut_2;
  reg        [7:0]    _26_9_inner_activation;
  reg        [7:0]    _26_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_9_inner_macOut;

  assign _zz__zz__26_9_inner_macOut = ($signed(io_mulInput) * $signed(_26_9_inner_activation));
  assign _zz__zz__26_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_9_inner_macOut)) ? 16'h007f : _zz__26_9_inner_macOut_2);
  assign _zz__26_9_inner_macOut_2 = (($signed(_zz__26_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_9_inner_activation;
    end else begin
      io_macOut = _26_9_inner_macOut;
    end
  end

  assign _zz__26_9_inner_macOut = ($signed(_zz__zz__26_9_inner_macOut) + $signed(_zz__zz__26_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_9_inner_activation <= 8'h00;
      _26_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_9_inner_activation <= io_addInput;
      end else begin
        _26_9_inner_macOut <= _zz__26_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_840 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_8_inner_macOut;
  wire       [15:0]   _zz__zz__26_8_inner_macOut_1;
  wire       [15:0]   _zz__26_8_inner_macOut_1;
  wire       [15:0]   _zz__26_8_inner_macOut_2;
  reg        [7:0]    _26_8_inner_activation;
  reg        [7:0]    _26_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_8_inner_macOut;

  assign _zz__zz__26_8_inner_macOut = ($signed(io_mulInput) * $signed(_26_8_inner_activation));
  assign _zz__zz__26_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_8_inner_macOut)) ? 16'h007f : _zz__26_8_inner_macOut_2);
  assign _zz__26_8_inner_macOut_2 = (($signed(_zz__26_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_8_inner_activation;
    end else begin
      io_macOut = _26_8_inner_macOut;
    end
  end

  assign _zz__26_8_inner_macOut = ($signed(_zz__zz__26_8_inner_macOut) + $signed(_zz__zz__26_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_8_inner_activation <= 8'h00;
      _26_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_8_inner_activation <= io_addInput;
      end else begin
        _26_8_inner_macOut <= _zz__26_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_839 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_7_inner_macOut;
  wire       [15:0]   _zz__zz__26_7_inner_macOut_1;
  wire       [15:0]   _zz__26_7_inner_macOut_1;
  wire       [15:0]   _zz__26_7_inner_macOut_2;
  reg        [7:0]    _26_7_inner_activation;
  reg        [7:0]    _26_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_7_inner_macOut;

  assign _zz__zz__26_7_inner_macOut = ($signed(io_mulInput) * $signed(_26_7_inner_activation));
  assign _zz__zz__26_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_7_inner_macOut)) ? 16'h007f : _zz__26_7_inner_macOut_2);
  assign _zz__26_7_inner_macOut_2 = (($signed(_zz__26_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_7_inner_activation;
    end else begin
      io_macOut = _26_7_inner_macOut;
    end
  end

  assign _zz__26_7_inner_macOut = ($signed(_zz__zz__26_7_inner_macOut) + $signed(_zz__zz__26_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_7_inner_activation <= 8'h00;
      _26_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_7_inner_activation <= io_addInput;
      end else begin
        _26_7_inner_macOut <= _zz__26_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_838 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_6_inner_macOut;
  wire       [15:0]   _zz__zz__26_6_inner_macOut_1;
  wire       [15:0]   _zz__26_6_inner_macOut_1;
  wire       [15:0]   _zz__26_6_inner_macOut_2;
  reg        [7:0]    _26_6_inner_activation;
  reg        [7:0]    _26_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_6_inner_macOut;

  assign _zz__zz__26_6_inner_macOut = ($signed(io_mulInput) * $signed(_26_6_inner_activation));
  assign _zz__zz__26_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_6_inner_macOut)) ? 16'h007f : _zz__26_6_inner_macOut_2);
  assign _zz__26_6_inner_macOut_2 = (($signed(_zz__26_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_6_inner_activation;
    end else begin
      io_macOut = _26_6_inner_macOut;
    end
  end

  assign _zz__26_6_inner_macOut = ($signed(_zz__zz__26_6_inner_macOut) + $signed(_zz__zz__26_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_6_inner_activation <= 8'h00;
      _26_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_6_inner_activation <= io_addInput;
      end else begin
        _26_6_inner_macOut <= _zz__26_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_837 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_5_inner_macOut;
  wire       [15:0]   _zz__zz__26_5_inner_macOut_1;
  wire       [15:0]   _zz__26_5_inner_macOut_1;
  wire       [15:0]   _zz__26_5_inner_macOut_2;
  reg        [7:0]    _26_5_inner_activation;
  reg        [7:0]    _26_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_5_inner_macOut;

  assign _zz__zz__26_5_inner_macOut = ($signed(io_mulInput) * $signed(_26_5_inner_activation));
  assign _zz__zz__26_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_5_inner_macOut)) ? 16'h007f : _zz__26_5_inner_macOut_2);
  assign _zz__26_5_inner_macOut_2 = (($signed(_zz__26_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_5_inner_activation;
    end else begin
      io_macOut = _26_5_inner_macOut;
    end
  end

  assign _zz__26_5_inner_macOut = ($signed(_zz__zz__26_5_inner_macOut) + $signed(_zz__zz__26_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_5_inner_activation <= 8'h00;
      _26_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_5_inner_activation <= io_addInput;
      end else begin
        _26_5_inner_macOut <= _zz__26_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_836 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_4_inner_macOut;
  wire       [15:0]   _zz__zz__26_4_inner_macOut_1;
  wire       [15:0]   _zz__26_4_inner_macOut_1;
  wire       [15:0]   _zz__26_4_inner_macOut_2;
  reg        [7:0]    _26_4_inner_activation;
  reg        [7:0]    _26_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_4_inner_macOut;

  assign _zz__zz__26_4_inner_macOut = ($signed(io_mulInput) * $signed(_26_4_inner_activation));
  assign _zz__zz__26_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_4_inner_macOut)) ? 16'h007f : _zz__26_4_inner_macOut_2);
  assign _zz__26_4_inner_macOut_2 = (($signed(_zz__26_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_4_inner_activation;
    end else begin
      io_macOut = _26_4_inner_macOut;
    end
  end

  assign _zz__26_4_inner_macOut = ($signed(_zz__zz__26_4_inner_macOut) + $signed(_zz__zz__26_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_4_inner_activation <= 8'h00;
      _26_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_4_inner_activation <= io_addInput;
      end else begin
        _26_4_inner_macOut <= _zz__26_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_835 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_3_inner_macOut;
  wire       [15:0]   _zz__zz__26_3_inner_macOut_1;
  wire       [15:0]   _zz__26_3_inner_macOut_1;
  wire       [15:0]   _zz__26_3_inner_macOut_2;
  reg        [7:0]    _26_3_inner_activation;
  reg        [7:0]    _26_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_3_inner_macOut;

  assign _zz__zz__26_3_inner_macOut = ($signed(io_mulInput) * $signed(_26_3_inner_activation));
  assign _zz__zz__26_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_3_inner_macOut)) ? 16'h007f : _zz__26_3_inner_macOut_2);
  assign _zz__26_3_inner_macOut_2 = (($signed(_zz__26_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_3_inner_activation;
    end else begin
      io_macOut = _26_3_inner_macOut;
    end
  end

  assign _zz__26_3_inner_macOut = ($signed(_zz__zz__26_3_inner_macOut) + $signed(_zz__zz__26_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_3_inner_activation <= 8'h00;
      _26_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_3_inner_activation <= io_addInput;
      end else begin
        _26_3_inner_macOut <= _zz__26_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_834 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_2_inner_macOut;
  wire       [15:0]   _zz__zz__26_2_inner_macOut_1;
  wire       [15:0]   _zz__26_2_inner_macOut_1;
  wire       [15:0]   _zz__26_2_inner_macOut_2;
  reg        [7:0]    _26_2_inner_activation;
  reg        [7:0]    _26_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_2_inner_macOut;

  assign _zz__zz__26_2_inner_macOut = ($signed(io_mulInput) * $signed(_26_2_inner_activation));
  assign _zz__zz__26_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_2_inner_macOut)) ? 16'h007f : _zz__26_2_inner_macOut_2);
  assign _zz__26_2_inner_macOut_2 = (($signed(_zz__26_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_2_inner_activation;
    end else begin
      io_macOut = _26_2_inner_macOut;
    end
  end

  assign _zz__26_2_inner_macOut = ($signed(_zz__zz__26_2_inner_macOut) + $signed(_zz__zz__26_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_2_inner_activation <= 8'h00;
      _26_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_2_inner_activation <= io_addInput;
      end else begin
        _26_2_inner_macOut <= _zz__26_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_833 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_1_inner_macOut;
  wire       [15:0]   _zz__zz__26_1_inner_macOut_1;
  wire       [15:0]   _zz__26_1_inner_macOut_1;
  wire       [15:0]   _zz__26_1_inner_macOut_2;
  reg        [7:0]    _26_1_inner_activation;
  reg        [7:0]    _26_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_1_inner_macOut;

  assign _zz__zz__26_1_inner_macOut = ($signed(io_mulInput) * $signed(_26_1_inner_activation));
  assign _zz__zz__26_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_1_inner_macOut)) ? 16'h007f : _zz__26_1_inner_macOut_2);
  assign _zz__26_1_inner_macOut_2 = (($signed(_zz__26_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_1_inner_activation;
    end else begin
      io_macOut = _26_1_inner_macOut;
    end
  end

  assign _zz__26_1_inner_macOut = ($signed(_zz__zz__26_1_inner_macOut) + $signed(_zz__zz__26_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_1_inner_activation <= 8'h00;
      _26_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_1_inner_activation <= io_addInput;
      end else begin
        _26_1_inner_macOut <= _zz__26_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_832 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__26_0_inner_macOut;
  wire       [15:0]   _zz__zz__26_0_inner_macOut_1;
  wire       [15:0]   _zz__26_0_inner_macOut_1;
  wire       [15:0]   _zz__26_0_inner_macOut_2;
  reg        [7:0]    _26_0_inner_activation;
  reg        [7:0]    _26_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__26_0_inner_macOut;

  assign _zz__zz__26_0_inner_macOut = ($signed(io_mulInput) * $signed(_26_0_inner_activation));
  assign _zz__zz__26_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__26_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__26_0_inner_macOut)) ? 16'h007f : _zz__26_0_inner_macOut_2);
  assign _zz__26_0_inner_macOut_2 = (($signed(_zz__26_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__26_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _26_0_inner_activation;
    end else begin
      io_macOut = _26_0_inner_macOut;
    end
  end

  assign _zz__26_0_inner_macOut = ($signed(_zz__zz__26_0_inner_macOut) + $signed(_zz__zz__26_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _26_0_inner_activation <= 8'h00;
      _26_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _26_0_inner_activation <= io_addInput;
      end else begin
        _26_0_inner_macOut <= _zz__26_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_831 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_31_inner_macOut;
  wire       [15:0]   _zz__zz__25_31_inner_macOut_1;
  wire       [15:0]   _zz__25_31_inner_macOut_1;
  wire       [15:0]   _zz__25_31_inner_macOut_2;
  reg        [7:0]    _25_31_inner_activation;
  reg        [7:0]    _25_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_31_inner_macOut;

  assign _zz__zz__25_31_inner_macOut = ($signed(io_mulInput) * $signed(_25_31_inner_activation));
  assign _zz__zz__25_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_31_inner_macOut)) ? 16'h007f : _zz__25_31_inner_macOut_2);
  assign _zz__25_31_inner_macOut_2 = (($signed(_zz__25_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_31_inner_activation;
    end else begin
      io_macOut = _25_31_inner_macOut;
    end
  end

  assign _zz__25_31_inner_macOut = ($signed(_zz__zz__25_31_inner_macOut) + $signed(_zz__zz__25_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_31_inner_activation <= 8'h00;
      _25_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_31_inner_activation <= io_addInput;
      end else begin
        _25_31_inner_macOut <= _zz__25_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_830 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_30_inner_macOut;
  wire       [15:0]   _zz__zz__25_30_inner_macOut_1;
  wire       [15:0]   _zz__25_30_inner_macOut_1;
  wire       [15:0]   _zz__25_30_inner_macOut_2;
  reg        [7:0]    _25_30_inner_activation;
  reg        [7:0]    _25_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_30_inner_macOut;

  assign _zz__zz__25_30_inner_macOut = ($signed(io_mulInput) * $signed(_25_30_inner_activation));
  assign _zz__zz__25_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_30_inner_macOut)) ? 16'h007f : _zz__25_30_inner_macOut_2);
  assign _zz__25_30_inner_macOut_2 = (($signed(_zz__25_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_30_inner_activation;
    end else begin
      io_macOut = _25_30_inner_macOut;
    end
  end

  assign _zz__25_30_inner_macOut = ($signed(_zz__zz__25_30_inner_macOut) + $signed(_zz__zz__25_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_30_inner_activation <= 8'h00;
      _25_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_30_inner_activation <= io_addInput;
      end else begin
        _25_30_inner_macOut <= _zz__25_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_829 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_29_inner_macOut;
  wire       [15:0]   _zz__zz__25_29_inner_macOut_1;
  wire       [15:0]   _zz__25_29_inner_macOut_1;
  wire       [15:0]   _zz__25_29_inner_macOut_2;
  reg        [7:0]    _25_29_inner_activation;
  reg        [7:0]    _25_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_29_inner_macOut;

  assign _zz__zz__25_29_inner_macOut = ($signed(io_mulInput) * $signed(_25_29_inner_activation));
  assign _zz__zz__25_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_29_inner_macOut)) ? 16'h007f : _zz__25_29_inner_macOut_2);
  assign _zz__25_29_inner_macOut_2 = (($signed(_zz__25_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_29_inner_activation;
    end else begin
      io_macOut = _25_29_inner_macOut;
    end
  end

  assign _zz__25_29_inner_macOut = ($signed(_zz__zz__25_29_inner_macOut) + $signed(_zz__zz__25_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_29_inner_activation <= 8'h00;
      _25_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_29_inner_activation <= io_addInput;
      end else begin
        _25_29_inner_macOut <= _zz__25_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_828 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_28_inner_macOut;
  wire       [15:0]   _zz__zz__25_28_inner_macOut_1;
  wire       [15:0]   _zz__25_28_inner_macOut_1;
  wire       [15:0]   _zz__25_28_inner_macOut_2;
  reg        [7:0]    _25_28_inner_activation;
  reg        [7:0]    _25_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_28_inner_macOut;

  assign _zz__zz__25_28_inner_macOut = ($signed(io_mulInput) * $signed(_25_28_inner_activation));
  assign _zz__zz__25_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_28_inner_macOut)) ? 16'h007f : _zz__25_28_inner_macOut_2);
  assign _zz__25_28_inner_macOut_2 = (($signed(_zz__25_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_28_inner_activation;
    end else begin
      io_macOut = _25_28_inner_macOut;
    end
  end

  assign _zz__25_28_inner_macOut = ($signed(_zz__zz__25_28_inner_macOut) + $signed(_zz__zz__25_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_28_inner_activation <= 8'h00;
      _25_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_28_inner_activation <= io_addInput;
      end else begin
        _25_28_inner_macOut <= _zz__25_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_827 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_27_inner_macOut;
  wire       [15:0]   _zz__zz__25_27_inner_macOut_1;
  wire       [15:0]   _zz__25_27_inner_macOut_1;
  wire       [15:0]   _zz__25_27_inner_macOut_2;
  reg        [7:0]    _25_27_inner_activation;
  reg        [7:0]    _25_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_27_inner_macOut;

  assign _zz__zz__25_27_inner_macOut = ($signed(io_mulInput) * $signed(_25_27_inner_activation));
  assign _zz__zz__25_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_27_inner_macOut)) ? 16'h007f : _zz__25_27_inner_macOut_2);
  assign _zz__25_27_inner_macOut_2 = (($signed(_zz__25_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_27_inner_activation;
    end else begin
      io_macOut = _25_27_inner_macOut;
    end
  end

  assign _zz__25_27_inner_macOut = ($signed(_zz__zz__25_27_inner_macOut) + $signed(_zz__zz__25_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_27_inner_activation <= 8'h00;
      _25_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_27_inner_activation <= io_addInput;
      end else begin
        _25_27_inner_macOut <= _zz__25_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_826 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_26_inner_macOut;
  wire       [15:0]   _zz__zz__25_26_inner_macOut_1;
  wire       [15:0]   _zz__25_26_inner_macOut_1;
  wire       [15:0]   _zz__25_26_inner_macOut_2;
  reg        [7:0]    _25_26_inner_activation;
  reg        [7:0]    _25_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_26_inner_macOut;

  assign _zz__zz__25_26_inner_macOut = ($signed(io_mulInput) * $signed(_25_26_inner_activation));
  assign _zz__zz__25_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_26_inner_macOut)) ? 16'h007f : _zz__25_26_inner_macOut_2);
  assign _zz__25_26_inner_macOut_2 = (($signed(_zz__25_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_26_inner_activation;
    end else begin
      io_macOut = _25_26_inner_macOut;
    end
  end

  assign _zz__25_26_inner_macOut = ($signed(_zz__zz__25_26_inner_macOut) + $signed(_zz__zz__25_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_26_inner_activation <= 8'h00;
      _25_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_26_inner_activation <= io_addInput;
      end else begin
        _25_26_inner_macOut <= _zz__25_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_825 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_25_inner_macOut;
  wire       [15:0]   _zz__zz__25_25_inner_macOut_1;
  wire       [15:0]   _zz__25_25_inner_macOut_1;
  wire       [15:0]   _zz__25_25_inner_macOut_2;
  reg        [7:0]    _25_25_inner_activation;
  reg        [7:0]    _25_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_25_inner_macOut;

  assign _zz__zz__25_25_inner_macOut = ($signed(io_mulInput) * $signed(_25_25_inner_activation));
  assign _zz__zz__25_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_25_inner_macOut)) ? 16'h007f : _zz__25_25_inner_macOut_2);
  assign _zz__25_25_inner_macOut_2 = (($signed(_zz__25_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_25_inner_activation;
    end else begin
      io_macOut = _25_25_inner_macOut;
    end
  end

  assign _zz__25_25_inner_macOut = ($signed(_zz__zz__25_25_inner_macOut) + $signed(_zz__zz__25_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_25_inner_activation <= 8'h00;
      _25_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_25_inner_activation <= io_addInput;
      end else begin
        _25_25_inner_macOut <= _zz__25_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_824 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_24_inner_macOut;
  wire       [15:0]   _zz__zz__25_24_inner_macOut_1;
  wire       [15:0]   _zz__25_24_inner_macOut_1;
  wire       [15:0]   _zz__25_24_inner_macOut_2;
  reg        [7:0]    _25_24_inner_activation;
  reg        [7:0]    _25_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_24_inner_macOut;

  assign _zz__zz__25_24_inner_macOut = ($signed(io_mulInput) * $signed(_25_24_inner_activation));
  assign _zz__zz__25_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_24_inner_macOut)) ? 16'h007f : _zz__25_24_inner_macOut_2);
  assign _zz__25_24_inner_macOut_2 = (($signed(_zz__25_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_24_inner_activation;
    end else begin
      io_macOut = _25_24_inner_macOut;
    end
  end

  assign _zz__25_24_inner_macOut = ($signed(_zz__zz__25_24_inner_macOut) + $signed(_zz__zz__25_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_24_inner_activation <= 8'h00;
      _25_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_24_inner_activation <= io_addInput;
      end else begin
        _25_24_inner_macOut <= _zz__25_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_823 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_23_inner_macOut;
  wire       [15:0]   _zz__zz__25_23_inner_macOut_1;
  wire       [15:0]   _zz__25_23_inner_macOut_1;
  wire       [15:0]   _zz__25_23_inner_macOut_2;
  reg        [7:0]    _25_23_inner_activation;
  reg        [7:0]    _25_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_23_inner_macOut;

  assign _zz__zz__25_23_inner_macOut = ($signed(io_mulInput) * $signed(_25_23_inner_activation));
  assign _zz__zz__25_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_23_inner_macOut)) ? 16'h007f : _zz__25_23_inner_macOut_2);
  assign _zz__25_23_inner_macOut_2 = (($signed(_zz__25_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_23_inner_activation;
    end else begin
      io_macOut = _25_23_inner_macOut;
    end
  end

  assign _zz__25_23_inner_macOut = ($signed(_zz__zz__25_23_inner_macOut) + $signed(_zz__zz__25_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_23_inner_activation <= 8'h00;
      _25_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_23_inner_activation <= io_addInput;
      end else begin
        _25_23_inner_macOut <= _zz__25_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_822 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_22_inner_macOut;
  wire       [15:0]   _zz__zz__25_22_inner_macOut_1;
  wire       [15:0]   _zz__25_22_inner_macOut_1;
  wire       [15:0]   _zz__25_22_inner_macOut_2;
  reg        [7:0]    _25_22_inner_activation;
  reg        [7:0]    _25_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_22_inner_macOut;

  assign _zz__zz__25_22_inner_macOut = ($signed(io_mulInput) * $signed(_25_22_inner_activation));
  assign _zz__zz__25_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_22_inner_macOut)) ? 16'h007f : _zz__25_22_inner_macOut_2);
  assign _zz__25_22_inner_macOut_2 = (($signed(_zz__25_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_22_inner_activation;
    end else begin
      io_macOut = _25_22_inner_macOut;
    end
  end

  assign _zz__25_22_inner_macOut = ($signed(_zz__zz__25_22_inner_macOut) + $signed(_zz__zz__25_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_22_inner_activation <= 8'h00;
      _25_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_22_inner_activation <= io_addInput;
      end else begin
        _25_22_inner_macOut <= _zz__25_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_821 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_21_inner_macOut;
  wire       [15:0]   _zz__zz__25_21_inner_macOut_1;
  wire       [15:0]   _zz__25_21_inner_macOut_1;
  wire       [15:0]   _zz__25_21_inner_macOut_2;
  reg        [7:0]    _25_21_inner_activation;
  reg        [7:0]    _25_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_21_inner_macOut;

  assign _zz__zz__25_21_inner_macOut = ($signed(io_mulInput) * $signed(_25_21_inner_activation));
  assign _zz__zz__25_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_21_inner_macOut)) ? 16'h007f : _zz__25_21_inner_macOut_2);
  assign _zz__25_21_inner_macOut_2 = (($signed(_zz__25_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_21_inner_activation;
    end else begin
      io_macOut = _25_21_inner_macOut;
    end
  end

  assign _zz__25_21_inner_macOut = ($signed(_zz__zz__25_21_inner_macOut) + $signed(_zz__zz__25_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_21_inner_activation <= 8'h00;
      _25_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_21_inner_activation <= io_addInput;
      end else begin
        _25_21_inner_macOut <= _zz__25_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_820 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_20_inner_macOut;
  wire       [15:0]   _zz__zz__25_20_inner_macOut_1;
  wire       [15:0]   _zz__25_20_inner_macOut_1;
  wire       [15:0]   _zz__25_20_inner_macOut_2;
  reg        [7:0]    _25_20_inner_activation;
  reg        [7:0]    _25_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_20_inner_macOut;

  assign _zz__zz__25_20_inner_macOut = ($signed(io_mulInput) * $signed(_25_20_inner_activation));
  assign _zz__zz__25_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_20_inner_macOut)) ? 16'h007f : _zz__25_20_inner_macOut_2);
  assign _zz__25_20_inner_macOut_2 = (($signed(_zz__25_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_20_inner_activation;
    end else begin
      io_macOut = _25_20_inner_macOut;
    end
  end

  assign _zz__25_20_inner_macOut = ($signed(_zz__zz__25_20_inner_macOut) + $signed(_zz__zz__25_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_20_inner_activation <= 8'h00;
      _25_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_20_inner_activation <= io_addInput;
      end else begin
        _25_20_inner_macOut <= _zz__25_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_819 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_19_inner_macOut;
  wire       [15:0]   _zz__zz__25_19_inner_macOut_1;
  wire       [15:0]   _zz__25_19_inner_macOut_1;
  wire       [15:0]   _zz__25_19_inner_macOut_2;
  reg        [7:0]    _25_19_inner_activation;
  reg        [7:0]    _25_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_19_inner_macOut;

  assign _zz__zz__25_19_inner_macOut = ($signed(io_mulInput) * $signed(_25_19_inner_activation));
  assign _zz__zz__25_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_19_inner_macOut)) ? 16'h007f : _zz__25_19_inner_macOut_2);
  assign _zz__25_19_inner_macOut_2 = (($signed(_zz__25_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_19_inner_activation;
    end else begin
      io_macOut = _25_19_inner_macOut;
    end
  end

  assign _zz__25_19_inner_macOut = ($signed(_zz__zz__25_19_inner_macOut) + $signed(_zz__zz__25_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_19_inner_activation <= 8'h00;
      _25_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_19_inner_activation <= io_addInput;
      end else begin
        _25_19_inner_macOut <= _zz__25_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_818 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_18_inner_macOut;
  wire       [15:0]   _zz__zz__25_18_inner_macOut_1;
  wire       [15:0]   _zz__25_18_inner_macOut_1;
  wire       [15:0]   _zz__25_18_inner_macOut_2;
  reg        [7:0]    _25_18_inner_activation;
  reg        [7:0]    _25_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_18_inner_macOut;

  assign _zz__zz__25_18_inner_macOut = ($signed(io_mulInput) * $signed(_25_18_inner_activation));
  assign _zz__zz__25_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_18_inner_macOut)) ? 16'h007f : _zz__25_18_inner_macOut_2);
  assign _zz__25_18_inner_macOut_2 = (($signed(_zz__25_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_18_inner_activation;
    end else begin
      io_macOut = _25_18_inner_macOut;
    end
  end

  assign _zz__25_18_inner_macOut = ($signed(_zz__zz__25_18_inner_macOut) + $signed(_zz__zz__25_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_18_inner_activation <= 8'h00;
      _25_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_18_inner_activation <= io_addInput;
      end else begin
        _25_18_inner_macOut <= _zz__25_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_817 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_17_inner_macOut;
  wire       [15:0]   _zz__zz__25_17_inner_macOut_1;
  wire       [15:0]   _zz__25_17_inner_macOut_1;
  wire       [15:0]   _zz__25_17_inner_macOut_2;
  reg        [7:0]    _25_17_inner_activation;
  reg        [7:0]    _25_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_17_inner_macOut;

  assign _zz__zz__25_17_inner_macOut = ($signed(io_mulInput) * $signed(_25_17_inner_activation));
  assign _zz__zz__25_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_17_inner_macOut)) ? 16'h007f : _zz__25_17_inner_macOut_2);
  assign _zz__25_17_inner_macOut_2 = (($signed(_zz__25_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_17_inner_activation;
    end else begin
      io_macOut = _25_17_inner_macOut;
    end
  end

  assign _zz__25_17_inner_macOut = ($signed(_zz__zz__25_17_inner_macOut) + $signed(_zz__zz__25_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_17_inner_activation <= 8'h00;
      _25_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_17_inner_activation <= io_addInput;
      end else begin
        _25_17_inner_macOut <= _zz__25_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_816 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_16_inner_macOut;
  wire       [15:0]   _zz__zz__25_16_inner_macOut_1;
  wire       [15:0]   _zz__25_16_inner_macOut_1;
  wire       [15:0]   _zz__25_16_inner_macOut_2;
  reg        [7:0]    _25_16_inner_activation;
  reg        [7:0]    _25_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_16_inner_macOut;

  assign _zz__zz__25_16_inner_macOut = ($signed(io_mulInput) * $signed(_25_16_inner_activation));
  assign _zz__zz__25_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_16_inner_macOut)) ? 16'h007f : _zz__25_16_inner_macOut_2);
  assign _zz__25_16_inner_macOut_2 = (($signed(_zz__25_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_16_inner_activation;
    end else begin
      io_macOut = _25_16_inner_macOut;
    end
  end

  assign _zz__25_16_inner_macOut = ($signed(_zz__zz__25_16_inner_macOut) + $signed(_zz__zz__25_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_16_inner_activation <= 8'h00;
      _25_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_16_inner_activation <= io_addInput;
      end else begin
        _25_16_inner_macOut <= _zz__25_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_815 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_15_inner_macOut;
  wire       [15:0]   _zz__zz__25_15_inner_macOut_1;
  wire       [15:0]   _zz__25_15_inner_macOut_1;
  wire       [15:0]   _zz__25_15_inner_macOut_2;
  reg        [7:0]    _25_15_inner_activation;
  reg        [7:0]    _25_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_15_inner_macOut;

  assign _zz__zz__25_15_inner_macOut = ($signed(io_mulInput) * $signed(_25_15_inner_activation));
  assign _zz__zz__25_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_15_inner_macOut)) ? 16'h007f : _zz__25_15_inner_macOut_2);
  assign _zz__25_15_inner_macOut_2 = (($signed(_zz__25_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_15_inner_activation;
    end else begin
      io_macOut = _25_15_inner_macOut;
    end
  end

  assign _zz__25_15_inner_macOut = ($signed(_zz__zz__25_15_inner_macOut) + $signed(_zz__zz__25_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_15_inner_activation <= 8'h00;
      _25_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_15_inner_activation <= io_addInput;
      end else begin
        _25_15_inner_macOut <= _zz__25_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_814 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_14_inner_macOut;
  wire       [15:0]   _zz__zz__25_14_inner_macOut_1;
  wire       [15:0]   _zz__25_14_inner_macOut_1;
  wire       [15:0]   _zz__25_14_inner_macOut_2;
  reg        [7:0]    _25_14_inner_activation;
  reg        [7:0]    _25_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_14_inner_macOut;

  assign _zz__zz__25_14_inner_macOut = ($signed(io_mulInput) * $signed(_25_14_inner_activation));
  assign _zz__zz__25_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_14_inner_macOut)) ? 16'h007f : _zz__25_14_inner_macOut_2);
  assign _zz__25_14_inner_macOut_2 = (($signed(_zz__25_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_14_inner_activation;
    end else begin
      io_macOut = _25_14_inner_macOut;
    end
  end

  assign _zz__25_14_inner_macOut = ($signed(_zz__zz__25_14_inner_macOut) + $signed(_zz__zz__25_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_14_inner_activation <= 8'h00;
      _25_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_14_inner_activation <= io_addInput;
      end else begin
        _25_14_inner_macOut <= _zz__25_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_813 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_13_inner_macOut;
  wire       [15:0]   _zz__zz__25_13_inner_macOut_1;
  wire       [15:0]   _zz__25_13_inner_macOut_1;
  wire       [15:0]   _zz__25_13_inner_macOut_2;
  reg        [7:0]    _25_13_inner_activation;
  reg        [7:0]    _25_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_13_inner_macOut;

  assign _zz__zz__25_13_inner_macOut = ($signed(io_mulInput) * $signed(_25_13_inner_activation));
  assign _zz__zz__25_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_13_inner_macOut)) ? 16'h007f : _zz__25_13_inner_macOut_2);
  assign _zz__25_13_inner_macOut_2 = (($signed(_zz__25_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_13_inner_activation;
    end else begin
      io_macOut = _25_13_inner_macOut;
    end
  end

  assign _zz__25_13_inner_macOut = ($signed(_zz__zz__25_13_inner_macOut) + $signed(_zz__zz__25_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_13_inner_activation <= 8'h00;
      _25_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_13_inner_activation <= io_addInput;
      end else begin
        _25_13_inner_macOut <= _zz__25_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_812 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_12_inner_macOut;
  wire       [15:0]   _zz__zz__25_12_inner_macOut_1;
  wire       [15:0]   _zz__25_12_inner_macOut_1;
  wire       [15:0]   _zz__25_12_inner_macOut_2;
  reg        [7:0]    _25_12_inner_activation;
  reg        [7:0]    _25_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_12_inner_macOut;

  assign _zz__zz__25_12_inner_macOut = ($signed(io_mulInput) * $signed(_25_12_inner_activation));
  assign _zz__zz__25_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_12_inner_macOut)) ? 16'h007f : _zz__25_12_inner_macOut_2);
  assign _zz__25_12_inner_macOut_2 = (($signed(_zz__25_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_12_inner_activation;
    end else begin
      io_macOut = _25_12_inner_macOut;
    end
  end

  assign _zz__25_12_inner_macOut = ($signed(_zz__zz__25_12_inner_macOut) + $signed(_zz__zz__25_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_12_inner_activation <= 8'h00;
      _25_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_12_inner_activation <= io_addInput;
      end else begin
        _25_12_inner_macOut <= _zz__25_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_811 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_11_inner_macOut;
  wire       [15:0]   _zz__zz__25_11_inner_macOut_1;
  wire       [15:0]   _zz__25_11_inner_macOut_1;
  wire       [15:0]   _zz__25_11_inner_macOut_2;
  reg        [7:0]    _25_11_inner_activation;
  reg        [7:0]    _25_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_11_inner_macOut;

  assign _zz__zz__25_11_inner_macOut = ($signed(io_mulInput) * $signed(_25_11_inner_activation));
  assign _zz__zz__25_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_11_inner_macOut)) ? 16'h007f : _zz__25_11_inner_macOut_2);
  assign _zz__25_11_inner_macOut_2 = (($signed(_zz__25_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_11_inner_activation;
    end else begin
      io_macOut = _25_11_inner_macOut;
    end
  end

  assign _zz__25_11_inner_macOut = ($signed(_zz__zz__25_11_inner_macOut) + $signed(_zz__zz__25_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_11_inner_activation <= 8'h00;
      _25_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_11_inner_activation <= io_addInput;
      end else begin
        _25_11_inner_macOut <= _zz__25_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_810 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_10_inner_macOut;
  wire       [15:0]   _zz__zz__25_10_inner_macOut_1;
  wire       [15:0]   _zz__25_10_inner_macOut_1;
  wire       [15:0]   _zz__25_10_inner_macOut_2;
  reg        [7:0]    _25_10_inner_activation;
  reg        [7:0]    _25_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_10_inner_macOut;

  assign _zz__zz__25_10_inner_macOut = ($signed(io_mulInput) * $signed(_25_10_inner_activation));
  assign _zz__zz__25_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_10_inner_macOut)) ? 16'h007f : _zz__25_10_inner_macOut_2);
  assign _zz__25_10_inner_macOut_2 = (($signed(_zz__25_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_10_inner_activation;
    end else begin
      io_macOut = _25_10_inner_macOut;
    end
  end

  assign _zz__25_10_inner_macOut = ($signed(_zz__zz__25_10_inner_macOut) + $signed(_zz__zz__25_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_10_inner_activation <= 8'h00;
      _25_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_10_inner_activation <= io_addInput;
      end else begin
        _25_10_inner_macOut <= _zz__25_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_809 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_9_inner_macOut;
  wire       [15:0]   _zz__zz__25_9_inner_macOut_1;
  wire       [15:0]   _zz__25_9_inner_macOut_1;
  wire       [15:0]   _zz__25_9_inner_macOut_2;
  reg        [7:0]    _25_9_inner_activation;
  reg        [7:0]    _25_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_9_inner_macOut;

  assign _zz__zz__25_9_inner_macOut = ($signed(io_mulInput) * $signed(_25_9_inner_activation));
  assign _zz__zz__25_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_9_inner_macOut)) ? 16'h007f : _zz__25_9_inner_macOut_2);
  assign _zz__25_9_inner_macOut_2 = (($signed(_zz__25_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_9_inner_activation;
    end else begin
      io_macOut = _25_9_inner_macOut;
    end
  end

  assign _zz__25_9_inner_macOut = ($signed(_zz__zz__25_9_inner_macOut) + $signed(_zz__zz__25_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_9_inner_activation <= 8'h00;
      _25_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_9_inner_activation <= io_addInput;
      end else begin
        _25_9_inner_macOut <= _zz__25_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_808 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_8_inner_macOut;
  wire       [15:0]   _zz__zz__25_8_inner_macOut_1;
  wire       [15:0]   _zz__25_8_inner_macOut_1;
  wire       [15:0]   _zz__25_8_inner_macOut_2;
  reg        [7:0]    _25_8_inner_activation;
  reg        [7:0]    _25_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_8_inner_macOut;

  assign _zz__zz__25_8_inner_macOut = ($signed(io_mulInput) * $signed(_25_8_inner_activation));
  assign _zz__zz__25_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_8_inner_macOut)) ? 16'h007f : _zz__25_8_inner_macOut_2);
  assign _zz__25_8_inner_macOut_2 = (($signed(_zz__25_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_8_inner_activation;
    end else begin
      io_macOut = _25_8_inner_macOut;
    end
  end

  assign _zz__25_8_inner_macOut = ($signed(_zz__zz__25_8_inner_macOut) + $signed(_zz__zz__25_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_8_inner_activation <= 8'h00;
      _25_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_8_inner_activation <= io_addInput;
      end else begin
        _25_8_inner_macOut <= _zz__25_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_807 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_7_inner_macOut;
  wire       [15:0]   _zz__zz__25_7_inner_macOut_1;
  wire       [15:0]   _zz__25_7_inner_macOut_1;
  wire       [15:0]   _zz__25_7_inner_macOut_2;
  reg        [7:0]    _25_7_inner_activation;
  reg        [7:0]    _25_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_7_inner_macOut;

  assign _zz__zz__25_7_inner_macOut = ($signed(io_mulInput) * $signed(_25_7_inner_activation));
  assign _zz__zz__25_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_7_inner_macOut)) ? 16'h007f : _zz__25_7_inner_macOut_2);
  assign _zz__25_7_inner_macOut_2 = (($signed(_zz__25_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_7_inner_activation;
    end else begin
      io_macOut = _25_7_inner_macOut;
    end
  end

  assign _zz__25_7_inner_macOut = ($signed(_zz__zz__25_7_inner_macOut) + $signed(_zz__zz__25_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_7_inner_activation <= 8'h00;
      _25_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_7_inner_activation <= io_addInput;
      end else begin
        _25_7_inner_macOut <= _zz__25_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_806 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_6_inner_macOut;
  wire       [15:0]   _zz__zz__25_6_inner_macOut_1;
  wire       [15:0]   _zz__25_6_inner_macOut_1;
  wire       [15:0]   _zz__25_6_inner_macOut_2;
  reg        [7:0]    _25_6_inner_activation;
  reg        [7:0]    _25_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_6_inner_macOut;

  assign _zz__zz__25_6_inner_macOut = ($signed(io_mulInput) * $signed(_25_6_inner_activation));
  assign _zz__zz__25_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_6_inner_macOut)) ? 16'h007f : _zz__25_6_inner_macOut_2);
  assign _zz__25_6_inner_macOut_2 = (($signed(_zz__25_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_6_inner_activation;
    end else begin
      io_macOut = _25_6_inner_macOut;
    end
  end

  assign _zz__25_6_inner_macOut = ($signed(_zz__zz__25_6_inner_macOut) + $signed(_zz__zz__25_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_6_inner_activation <= 8'h00;
      _25_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_6_inner_activation <= io_addInput;
      end else begin
        _25_6_inner_macOut <= _zz__25_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_805 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_5_inner_macOut;
  wire       [15:0]   _zz__zz__25_5_inner_macOut_1;
  wire       [15:0]   _zz__25_5_inner_macOut_1;
  wire       [15:0]   _zz__25_5_inner_macOut_2;
  reg        [7:0]    _25_5_inner_activation;
  reg        [7:0]    _25_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_5_inner_macOut;

  assign _zz__zz__25_5_inner_macOut = ($signed(io_mulInput) * $signed(_25_5_inner_activation));
  assign _zz__zz__25_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_5_inner_macOut)) ? 16'h007f : _zz__25_5_inner_macOut_2);
  assign _zz__25_5_inner_macOut_2 = (($signed(_zz__25_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_5_inner_activation;
    end else begin
      io_macOut = _25_5_inner_macOut;
    end
  end

  assign _zz__25_5_inner_macOut = ($signed(_zz__zz__25_5_inner_macOut) + $signed(_zz__zz__25_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_5_inner_activation <= 8'h00;
      _25_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_5_inner_activation <= io_addInput;
      end else begin
        _25_5_inner_macOut <= _zz__25_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_804 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_4_inner_macOut;
  wire       [15:0]   _zz__zz__25_4_inner_macOut_1;
  wire       [15:0]   _zz__25_4_inner_macOut_1;
  wire       [15:0]   _zz__25_4_inner_macOut_2;
  reg        [7:0]    _25_4_inner_activation;
  reg        [7:0]    _25_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_4_inner_macOut;

  assign _zz__zz__25_4_inner_macOut = ($signed(io_mulInput) * $signed(_25_4_inner_activation));
  assign _zz__zz__25_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_4_inner_macOut)) ? 16'h007f : _zz__25_4_inner_macOut_2);
  assign _zz__25_4_inner_macOut_2 = (($signed(_zz__25_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_4_inner_activation;
    end else begin
      io_macOut = _25_4_inner_macOut;
    end
  end

  assign _zz__25_4_inner_macOut = ($signed(_zz__zz__25_4_inner_macOut) + $signed(_zz__zz__25_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_4_inner_activation <= 8'h00;
      _25_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_4_inner_activation <= io_addInput;
      end else begin
        _25_4_inner_macOut <= _zz__25_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_803 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_3_inner_macOut;
  wire       [15:0]   _zz__zz__25_3_inner_macOut_1;
  wire       [15:0]   _zz__25_3_inner_macOut_1;
  wire       [15:0]   _zz__25_3_inner_macOut_2;
  reg        [7:0]    _25_3_inner_activation;
  reg        [7:0]    _25_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_3_inner_macOut;

  assign _zz__zz__25_3_inner_macOut = ($signed(io_mulInput) * $signed(_25_3_inner_activation));
  assign _zz__zz__25_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_3_inner_macOut)) ? 16'h007f : _zz__25_3_inner_macOut_2);
  assign _zz__25_3_inner_macOut_2 = (($signed(_zz__25_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_3_inner_activation;
    end else begin
      io_macOut = _25_3_inner_macOut;
    end
  end

  assign _zz__25_3_inner_macOut = ($signed(_zz__zz__25_3_inner_macOut) + $signed(_zz__zz__25_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_3_inner_activation <= 8'h00;
      _25_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_3_inner_activation <= io_addInput;
      end else begin
        _25_3_inner_macOut <= _zz__25_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_802 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_2_inner_macOut;
  wire       [15:0]   _zz__zz__25_2_inner_macOut_1;
  wire       [15:0]   _zz__25_2_inner_macOut_1;
  wire       [15:0]   _zz__25_2_inner_macOut_2;
  reg        [7:0]    _25_2_inner_activation;
  reg        [7:0]    _25_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_2_inner_macOut;

  assign _zz__zz__25_2_inner_macOut = ($signed(io_mulInput) * $signed(_25_2_inner_activation));
  assign _zz__zz__25_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_2_inner_macOut)) ? 16'h007f : _zz__25_2_inner_macOut_2);
  assign _zz__25_2_inner_macOut_2 = (($signed(_zz__25_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_2_inner_activation;
    end else begin
      io_macOut = _25_2_inner_macOut;
    end
  end

  assign _zz__25_2_inner_macOut = ($signed(_zz__zz__25_2_inner_macOut) + $signed(_zz__zz__25_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_2_inner_activation <= 8'h00;
      _25_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_2_inner_activation <= io_addInput;
      end else begin
        _25_2_inner_macOut <= _zz__25_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_801 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_1_inner_macOut;
  wire       [15:0]   _zz__zz__25_1_inner_macOut_1;
  wire       [15:0]   _zz__25_1_inner_macOut_1;
  wire       [15:0]   _zz__25_1_inner_macOut_2;
  reg        [7:0]    _25_1_inner_activation;
  reg        [7:0]    _25_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_1_inner_macOut;

  assign _zz__zz__25_1_inner_macOut = ($signed(io_mulInput) * $signed(_25_1_inner_activation));
  assign _zz__zz__25_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_1_inner_macOut)) ? 16'h007f : _zz__25_1_inner_macOut_2);
  assign _zz__25_1_inner_macOut_2 = (($signed(_zz__25_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_1_inner_activation;
    end else begin
      io_macOut = _25_1_inner_macOut;
    end
  end

  assign _zz__25_1_inner_macOut = ($signed(_zz__zz__25_1_inner_macOut) + $signed(_zz__zz__25_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_1_inner_activation <= 8'h00;
      _25_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_1_inner_activation <= io_addInput;
      end else begin
        _25_1_inner_macOut <= _zz__25_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_800 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__25_0_inner_macOut;
  wire       [15:0]   _zz__zz__25_0_inner_macOut_1;
  wire       [15:0]   _zz__25_0_inner_macOut_1;
  wire       [15:0]   _zz__25_0_inner_macOut_2;
  reg        [7:0]    _25_0_inner_activation;
  reg        [7:0]    _25_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__25_0_inner_macOut;

  assign _zz__zz__25_0_inner_macOut = ($signed(io_mulInput) * $signed(_25_0_inner_activation));
  assign _zz__zz__25_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__25_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__25_0_inner_macOut)) ? 16'h007f : _zz__25_0_inner_macOut_2);
  assign _zz__25_0_inner_macOut_2 = (($signed(_zz__25_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__25_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _25_0_inner_activation;
    end else begin
      io_macOut = _25_0_inner_macOut;
    end
  end

  assign _zz__25_0_inner_macOut = ($signed(_zz__zz__25_0_inner_macOut) + $signed(_zz__zz__25_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _25_0_inner_activation <= 8'h00;
      _25_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _25_0_inner_activation <= io_addInput;
      end else begin
        _25_0_inner_macOut <= _zz__25_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_799 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_31_inner_macOut;
  wire       [15:0]   _zz__zz__24_31_inner_macOut_1;
  wire       [15:0]   _zz__24_31_inner_macOut_1;
  wire       [15:0]   _zz__24_31_inner_macOut_2;
  reg        [7:0]    _24_31_inner_activation;
  reg        [7:0]    _24_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_31_inner_macOut;

  assign _zz__zz__24_31_inner_macOut = ($signed(io_mulInput) * $signed(_24_31_inner_activation));
  assign _zz__zz__24_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_31_inner_macOut)) ? 16'h007f : _zz__24_31_inner_macOut_2);
  assign _zz__24_31_inner_macOut_2 = (($signed(_zz__24_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_31_inner_activation;
    end else begin
      io_macOut = _24_31_inner_macOut;
    end
  end

  assign _zz__24_31_inner_macOut = ($signed(_zz__zz__24_31_inner_macOut) + $signed(_zz__zz__24_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_31_inner_activation <= 8'h00;
      _24_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_31_inner_activation <= io_addInput;
      end else begin
        _24_31_inner_macOut <= _zz__24_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_798 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_30_inner_macOut;
  wire       [15:0]   _zz__zz__24_30_inner_macOut_1;
  wire       [15:0]   _zz__24_30_inner_macOut_1;
  wire       [15:0]   _zz__24_30_inner_macOut_2;
  reg        [7:0]    _24_30_inner_activation;
  reg        [7:0]    _24_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_30_inner_macOut;

  assign _zz__zz__24_30_inner_macOut = ($signed(io_mulInput) * $signed(_24_30_inner_activation));
  assign _zz__zz__24_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_30_inner_macOut)) ? 16'h007f : _zz__24_30_inner_macOut_2);
  assign _zz__24_30_inner_macOut_2 = (($signed(_zz__24_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_30_inner_activation;
    end else begin
      io_macOut = _24_30_inner_macOut;
    end
  end

  assign _zz__24_30_inner_macOut = ($signed(_zz__zz__24_30_inner_macOut) + $signed(_zz__zz__24_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_30_inner_activation <= 8'h00;
      _24_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_30_inner_activation <= io_addInput;
      end else begin
        _24_30_inner_macOut <= _zz__24_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_797 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_29_inner_macOut;
  wire       [15:0]   _zz__zz__24_29_inner_macOut_1;
  wire       [15:0]   _zz__24_29_inner_macOut_1;
  wire       [15:0]   _zz__24_29_inner_macOut_2;
  reg        [7:0]    _24_29_inner_activation;
  reg        [7:0]    _24_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_29_inner_macOut;

  assign _zz__zz__24_29_inner_macOut = ($signed(io_mulInput) * $signed(_24_29_inner_activation));
  assign _zz__zz__24_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_29_inner_macOut)) ? 16'h007f : _zz__24_29_inner_macOut_2);
  assign _zz__24_29_inner_macOut_2 = (($signed(_zz__24_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_29_inner_activation;
    end else begin
      io_macOut = _24_29_inner_macOut;
    end
  end

  assign _zz__24_29_inner_macOut = ($signed(_zz__zz__24_29_inner_macOut) + $signed(_zz__zz__24_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_29_inner_activation <= 8'h00;
      _24_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_29_inner_activation <= io_addInput;
      end else begin
        _24_29_inner_macOut <= _zz__24_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_796 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_28_inner_macOut;
  wire       [15:0]   _zz__zz__24_28_inner_macOut_1;
  wire       [15:0]   _zz__24_28_inner_macOut_1;
  wire       [15:0]   _zz__24_28_inner_macOut_2;
  reg        [7:0]    _24_28_inner_activation;
  reg        [7:0]    _24_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_28_inner_macOut;

  assign _zz__zz__24_28_inner_macOut = ($signed(io_mulInput) * $signed(_24_28_inner_activation));
  assign _zz__zz__24_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_28_inner_macOut)) ? 16'h007f : _zz__24_28_inner_macOut_2);
  assign _zz__24_28_inner_macOut_2 = (($signed(_zz__24_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_28_inner_activation;
    end else begin
      io_macOut = _24_28_inner_macOut;
    end
  end

  assign _zz__24_28_inner_macOut = ($signed(_zz__zz__24_28_inner_macOut) + $signed(_zz__zz__24_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_28_inner_activation <= 8'h00;
      _24_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_28_inner_activation <= io_addInput;
      end else begin
        _24_28_inner_macOut <= _zz__24_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_795 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_27_inner_macOut;
  wire       [15:0]   _zz__zz__24_27_inner_macOut_1;
  wire       [15:0]   _zz__24_27_inner_macOut_1;
  wire       [15:0]   _zz__24_27_inner_macOut_2;
  reg        [7:0]    _24_27_inner_activation;
  reg        [7:0]    _24_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_27_inner_macOut;

  assign _zz__zz__24_27_inner_macOut = ($signed(io_mulInput) * $signed(_24_27_inner_activation));
  assign _zz__zz__24_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_27_inner_macOut)) ? 16'h007f : _zz__24_27_inner_macOut_2);
  assign _zz__24_27_inner_macOut_2 = (($signed(_zz__24_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_27_inner_activation;
    end else begin
      io_macOut = _24_27_inner_macOut;
    end
  end

  assign _zz__24_27_inner_macOut = ($signed(_zz__zz__24_27_inner_macOut) + $signed(_zz__zz__24_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_27_inner_activation <= 8'h00;
      _24_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_27_inner_activation <= io_addInput;
      end else begin
        _24_27_inner_macOut <= _zz__24_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_794 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_26_inner_macOut;
  wire       [15:0]   _zz__zz__24_26_inner_macOut_1;
  wire       [15:0]   _zz__24_26_inner_macOut_1;
  wire       [15:0]   _zz__24_26_inner_macOut_2;
  reg        [7:0]    _24_26_inner_activation;
  reg        [7:0]    _24_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_26_inner_macOut;

  assign _zz__zz__24_26_inner_macOut = ($signed(io_mulInput) * $signed(_24_26_inner_activation));
  assign _zz__zz__24_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_26_inner_macOut)) ? 16'h007f : _zz__24_26_inner_macOut_2);
  assign _zz__24_26_inner_macOut_2 = (($signed(_zz__24_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_26_inner_activation;
    end else begin
      io_macOut = _24_26_inner_macOut;
    end
  end

  assign _zz__24_26_inner_macOut = ($signed(_zz__zz__24_26_inner_macOut) + $signed(_zz__zz__24_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_26_inner_activation <= 8'h00;
      _24_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_26_inner_activation <= io_addInput;
      end else begin
        _24_26_inner_macOut <= _zz__24_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_793 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_25_inner_macOut;
  wire       [15:0]   _zz__zz__24_25_inner_macOut_1;
  wire       [15:0]   _zz__24_25_inner_macOut_1;
  wire       [15:0]   _zz__24_25_inner_macOut_2;
  reg        [7:0]    _24_25_inner_activation;
  reg        [7:0]    _24_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_25_inner_macOut;

  assign _zz__zz__24_25_inner_macOut = ($signed(io_mulInput) * $signed(_24_25_inner_activation));
  assign _zz__zz__24_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_25_inner_macOut)) ? 16'h007f : _zz__24_25_inner_macOut_2);
  assign _zz__24_25_inner_macOut_2 = (($signed(_zz__24_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_25_inner_activation;
    end else begin
      io_macOut = _24_25_inner_macOut;
    end
  end

  assign _zz__24_25_inner_macOut = ($signed(_zz__zz__24_25_inner_macOut) + $signed(_zz__zz__24_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_25_inner_activation <= 8'h00;
      _24_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_25_inner_activation <= io_addInput;
      end else begin
        _24_25_inner_macOut <= _zz__24_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_792 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_24_inner_macOut;
  wire       [15:0]   _zz__zz__24_24_inner_macOut_1;
  wire       [15:0]   _zz__24_24_inner_macOut_1;
  wire       [15:0]   _zz__24_24_inner_macOut_2;
  reg        [7:0]    _24_24_inner_activation;
  reg        [7:0]    _24_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_24_inner_macOut;

  assign _zz__zz__24_24_inner_macOut = ($signed(io_mulInput) * $signed(_24_24_inner_activation));
  assign _zz__zz__24_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_24_inner_macOut)) ? 16'h007f : _zz__24_24_inner_macOut_2);
  assign _zz__24_24_inner_macOut_2 = (($signed(_zz__24_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_24_inner_activation;
    end else begin
      io_macOut = _24_24_inner_macOut;
    end
  end

  assign _zz__24_24_inner_macOut = ($signed(_zz__zz__24_24_inner_macOut) + $signed(_zz__zz__24_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_24_inner_activation <= 8'h00;
      _24_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_24_inner_activation <= io_addInput;
      end else begin
        _24_24_inner_macOut <= _zz__24_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_791 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_23_inner_macOut;
  wire       [15:0]   _zz__zz__24_23_inner_macOut_1;
  wire       [15:0]   _zz__24_23_inner_macOut_1;
  wire       [15:0]   _zz__24_23_inner_macOut_2;
  reg        [7:0]    _24_23_inner_activation;
  reg        [7:0]    _24_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_23_inner_macOut;

  assign _zz__zz__24_23_inner_macOut = ($signed(io_mulInput) * $signed(_24_23_inner_activation));
  assign _zz__zz__24_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_23_inner_macOut)) ? 16'h007f : _zz__24_23_inner_macOut_2);
  assign _zz__24_23_inner_macOut_2 = (($signed(_zz__24_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_23_inner_activation;
    end else begin
      io_macOut = _24_23_inner_macOut;
    end
  end

  assign _zz__24_23_inner_macOut = ($signed(_zz__zz__24_23_inner_macOut) + $signed(_zz__zz__24_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_23_inner_activation <= 8'h00;
      _24_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_23_inner_activation <= io_addInput;
      end else begin
        _24_23_inner_macOut <= _zz__24_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_790 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_22_inner_macOut;
  wire       [15:0]   _zz__zz__24_22_inner_macOut_1;
  wire       [15:0]   _zz__24_22_inner_macOut_1;
  wire       [15:0]   _zz__24_22_inner_macOut_2;
  reg        [7:0]    _24_22_inner_activation;
  reg        [7:0]    _24_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_22_inner_macOut;

  assign _zz__zz__24_22_inner_macOut = ($signed(io_mulInput) * $signed(_24_22_inner_activation));
  assign _zz__zz__24_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_22_inner_macOut)) ? 16'h007f : _zz__24_22_inner_macOut_2);
  assign _zz__24_22_inner_macOut_2 = (($signed(_zz__24_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_22_inner_activation;
    end else begin
      io_macOut = _24_22_inner_macOut;
    end
  end

  assign _zz__24_22_inner_macOut = ($signed(_zz__zz__24_22_inner_macOut) + $signed(_zz__zz__24_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_22_inner_activation <= 8'h00;
      _24_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_22_inner_activation <= io_addInput;
      end else begin
        _24_22_inner_macOut <= _zz__24_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_789 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_21_inner_macOut;
  wire       [15:0]   _zz__zz__24_21_inner_macOut_1;
  wire       [15:0]   _zz__24_21_inner_macOut_1;
  wire       [15:0]   _zz__24_21_inner_macOut_2;
  reg        [7:0]    _24_21_inner_activation;
  reg        [7:0]    _24_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_21_inner_macOut;

  assign _zz__zz__24_21_inner_macOut = ($signed(io_mulInput) * $signed(_24_21_inner_activation));
  assign _zz__zz__24_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_21_inner_macOut)) ? 16'h007f : _zz__24_21_inner_macOut_2);
  assign _zz__24_21_inner_macOut_2 = (($signed(_zz__24_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_21_inner_activation;
    end else begin
      io_macOut = _24_21_inner_macOut;
    end
  end

  assign _zz__24_21_inner_macOut = ($signed(_zz__zz__24_21_inner_macOut) + $signed(_zz__zz__24_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_21_inner_activation <= 8'h00;
      _24_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_21_inner_activation <= io_addInput;
      end else begin
        _24_21_inner_macOut <= _zz__24_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_788 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_20_inner_macOut;
  wire       [15:0]   _zz__zz__24_20_inner_macOut_1;
  wire       [15:0]   _zz__24_20_inner_macOut_1;
  wire       [15:0]   _zz__24_20_inner_macOut_2;
  reg        [7:0]    _24_20_inner_activation;
  reg        [7:0]    _24_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_20_inner_macOut;

  assign _zz__zz__24_20_inner_macOut = ($signed(io_mulInput) * $signed(_24_20_inner_activation));
  assign _zz__zz__24_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_20_inner_macOut)) ? 16'h007f : _zz__24_20_inner_macOut_2);
  assign _zz__24_20_inner_macOut_2 = (($signed(_zz__24_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_20_inner_activation;
    end else begin
      io_macOut = _24_20_inner_macOut;
    end
  end

  assign _zz__24_20_inner_macOut = ($signed(_zz__zz__24_20_inner_macOut) + $signed(_zz__zz__24_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_20_inner_activation <= 8'h00;
      _24_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_20_inner_activation <= io_addInput;
      end else begin
        _24_20_inner_macOut <= _zz__24_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_787 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_19_inner_macOut;
  wire       [15:0]   _zz__zz__24_19_inner_macOut_1;
  wire       [15:0]   _zz__24_19_inner_macOut_1;
  wire       [15:0]   _zz__24_19_inner_macOut_2;
  reg        [7:0]    _24_19_inner_activation;
  reg        [7:0]    _24_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_19_inner_macOut;

  assign _zz__zz__24_19_inner_macOut = ($signed(io_mulInput) * $signed(_24_19_inner_activation));
  assign _zz__zz__24_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_19_inner_macOut)) ? 16'h007f : _zz__24_19_inner_macOut_2);
  assign _zz__24_19_inner_macOut_2 = (($signed(_zz__24_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_19_inner_activation;
    end else begin
      io_macOut = _24_19_inner_macOut;
    end
  end

  assign _zz__24_19_inner_macOut = ($signed(_zz__zz__24_19_inner_macOut) + $signed(_zz__zz__24_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_19_inner_activation <= 8'h00;
      _24_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_19_inner_activation <= io_addInput;
      end else begin
        _24_19_inner_macOut <= _zz__24_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_786 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_18_inner_macOut;
  wire       [15:0]   _zz__zz__24_18_inner_macOut_1;
  wire       [15:0]   _zz__24_18_inner_macOut_1;
  wire       [15:0]   _zz__24_18_inner_macOut_2;
  reg        [7:0]    _24_18_inner_activation;
  reg        [7:0]    _24_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_18_inner_macOut;

  assign _zz__zz__24_18_inner_macOut = ($signed(io_mulInput) * $signed(_24_18_inner_activation));
  assign _zz__zz__24_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_18_inner_macOut)) ? 16'h007f : _zz__24_18_inner_macOut_2);
  assign _zz__24_18_inner_macOut_2 = (($signed(_zz__24_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_18_inner_activation;
    end else begin
      io_macOut = _24_18_inner_macOut;
    end
  end

  assign _zz__24_18_inner_macOut = ($signed(_zz__zz__24_18_inner_macOut) + $signed(_zz__zz__24_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_18_inner_activation <= 8'h00;
      _24_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_18_inner_activation <= io_addInput;
      end else begin
        _24_18_inner_macOut <= _zz__24_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_785 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_17_inner_macOut;
  wire       [15:0]   _zz__zz__24_17_inner_macOut_1;
  wire       [15:0]   _zz__24_17_inner_macOut_1;
  wire       [15:0]   _zz__24_17_inner_macOut_2;
  reg        [7:0]    _24_17_inner_activation;
  reg        [7:0]    _24_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_17_inner_macOut;

  assign _zz__zz__24_17_inner_macOut = ($signed(io_mulInput) * $signed(_24_17_inner_activation));
  assign _zz__zz__24_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_17_inner_macOut)) ? 16'h007f : _zz__24_17_inner_macOut_2);
  assign _zz__24_17_inner_macOut_2 = (($signed(_zz__24_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_17_inner_activation;
    end else begin
      io_macOut = _24_17_inner_macOut;
    end
  end

  assign _zz__24_17_inner_macOut = ($signed(_zz__zz__24_17_inner_macOut) + $signed(_zz__zz__24_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_17_inner_activation <= 8'h00;
      _24_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_17_inner_activation <= io_addInput;
      end else begin
        _24_17_inner_macOut <= _zz__24_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_784 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_16_inner_macOut;
  wire       [15:0]   _zz__zz__24_16_inner_macOut_1;
  wire       [15:0]   _zz__24_16_inner_macOut_1;
  wire       [15:0]   _zz__24_16_inner_macOut_2;
  reg        [7:0]    _24_16_inner_activation;
  reg        [7:0]    _24_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_16_inner_macOut;

  assign _zz__zz__24_16_inner_macOut = ($signed(io_mulInput) * $signed(_24_16_inner_activation));
  assign _zz__zz__24_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_16_inner_macOut)) ? 16'h007f : _zz__24_16_inner_macOut_2);
  assign _zz__24_16_inner_macOut_2 = (($signed(_zz__24_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_16_inner_activation;
    end else begin
      io_macOut = _24_16_inner_macOut;
    end
  end

  assign _zz__24_16_inner_macOut = ($signed(_zz__zz__24_16_inner_macOut) + $signed(_zz__zz__24_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_16_inner_activation <= 8'h00;
      _24_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_16_inner_activation <= io_addInput;
      end else begin
        _24_16_inner_macOut <= _zz__24_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_783 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_15_inner_macOut;
  wire       [15:0]   _zz__zz__24_15_inner_macOut_1;
  wire       [15:0]   _zz__24_15_inner_macOut_1;
  wire       [15:0]   _zz__24_15_inner_macOut_2;
  reg        [7:0]    _24_15_inner_activation;
  reg        [7:0]    _24_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_15_inner_macOut;

  assign _zz__zz__24_15_inner_macOut = ($signed(io_mulInput) * $signed(_24_15_inner_activation));
  assign _zz__zz__24_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_15_inner_macOut)) ? 16'h007f : _zz__24_15_inner_macOut_2);
  assign _zz__24_15_inner_macOut_2 = (($signed(_zz__24_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_15_inner_activation;
    end else begin
      io_macOut = _24_15_inner_macOut;
    end
  end

  assign _zz__24_15_inner_macOut = ($signed(_zz__zz__24_15_inner_macOut) + $signed(_zz__zz__24_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_15_inner_activation <= 8'h00;
      _24_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_15_inner_activation <= io_addInput;
      end else begin
        _24_15_inner_macOut <= _zz__24_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_782 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_14_inner_macOut;
  wire       [15:0]   _zz__zz__24_14_inner_macOut_1;
  wire       [15:0]   _zz__24_14_inner_macOut_1;
  wire       [15:0]   _zz__24_14_inner_macOut_2;
  reg        [7:0]    _24_14_inner_activation;
  reg        [7:0]    _24_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_14_inner_macOut;

  assign _zz__zz__24_14_inner_macOut = ($signed(io_mulInput) * $signed(_24_14_inner_activation));
  assign _zz__zz__24_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_14_inner_macOut)) ? 16'h007f : _zz__24_14_inner_macOut_2);
  assign _zz__24_14_inner_macOut_2 = (($signed(_zz__24_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_14_inner_activation;
    end else begin
      io_macOut = _24_14_inner_macOut;
    end
  end

  assign _zz__24_14_inner_macOut = ($signed(_zz__zz__24_14_inner_macOut) + $signed(_zz__zz__24_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_14_inner_activation <= 8'h00;
      _24_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_14_inner_activation <= io_addInput;
      end else begin
        _24_14_inner_macOut <= _zz__24_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_781 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_13_inner_macOut;
  wire       [15:0]   _zz__zz__24_13_inner_macOut_1;
  wire       [15:0]   _zz__24_13_inner_macOut_1;
  wire       [15:0]   _zz__24_13_inner_macOut_2;
  reg        [7:0]    _24_13_inner_activation;
  reg        [7:0]    _24_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_13_inner_macOut;

  assign _zz__zz__24_13_inner_macOut = ($signed(io_mulInput) * $signed(_24_13_inner_activation));
  assign _zz__zz__24_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_13_inner_macOut)) ? 16'h007f : _zz__24_13_inner_macOut_2);
  assign _zz__24_13_inner_macOut_2 = (($signed(_zz__24_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_13_inner_activation;
    end else begin
      io_macOut = _24_13_inner_macOut;
    end
  end

  assign _zz__24_13_inner_macOut = ($signed(_zz__zz__24_13_inner_macOut) + $signed(_zz__zz__24_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_13_inner_activation <= 8'h00;
      _24_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_13_inner_activation <= io_addInput;
      end else begin
        _24_13_inner_macOut <= _zz__24_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_780 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_12_inner_macOut;
  wire       [15:0]   _zz__zz__24_12_inner_macOut_1;
  wire       [15:0]   _zz__24_12_inner_macOut_1;
  wire       [15:0]   _zz__24_12_inner_macOut_2;
  reg        [7:0]    _24_12_inner_activation;
  reg        [7:0]    _24_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_12_inner_macOut;

  assign _zz__zz__24_12_inner_macOut = ($signed(io_mulInput) * $signed(_24_12_inner_activation));
  assign _zz__zz__24_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_12_inner_macOut)) ? 16'h007f : _zz__24_12_inner_macOut_2);
  assign _zz__24_12_inner_macOut_2 = (($signed(_zz__24_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_12_inner_activation;
    end else begin
      io_macOut = _24_12_inner_macOut;
    end
  end

  assign _zz__24_12_inner_macOut = ($signed(_zz__zz__24_12_inner_macOut) + $signed(_zz__zz__24_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_12_inner_activation <= 8'h00;
      _24_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_12_inner_activation <= io_addInput;
      end else begin
        _24_12_inner_macOut <= _zz__24_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_779 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_11_inner_macOut;
  wire       [15:0]   _zz__zz__24_11_inner_macOut_1;
  wire       [15:0]   _zz__24_11_inner_macOut_1;
  wire       [15:0]   _zz__24_11_inner_macOut_2;
  reg        [7:0]    _24_11_inner_activation;
  reg        [7:0]    _24_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_11_inner_macOut;

  assign _zz__zz__24_11_inner_macOut = ($signed(io_mulInput) * $signed(_24_11_inner_activation));
  assign _zz__zz__24_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_11_inner_macOut)) ? 16'h007f : _zz__24_11_inner_macOut_2);
  assign _zz__24_11_inner_macOut_2 = (($signed(_zz__24_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_11_inner_activation;
    end else begin
      io_macOut = _24_11_inner_macOut;
    end
  end

  assign _zz__24_11_inner_macOut = ($signed(_zz__zz__24_11_inner_macOut) + $signed(_zz__zz__24_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_11_inner_activation <= 8'h00;
      _24_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_11_inner_activation <= io_addInput;
      end else begin
        _24_11_inner_macOut <= _zz__24_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_778 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_10_inner_macOut;
  wire       [15:0]   _zz__zz__24_10_inner_macOut_1;
  wire       [15:0]   _zz__24_10_inner_macOut_1;
  wire       [15:0]   _zz__24_10_inner_macOut_2;
  reg        [7:0]    _24_10_inner_activation;
  reg        [7:0]    _24_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_10_inner_macOut;

  assign _zz__zz__24_10_inner_macOut = ($signed(io_mulInput) * $signed(_24_10_inner_activation));
  assign _zz__zz__24_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_10_inner_macOut)) ? 16'h007f : _zz__24_10_inner_macOut_2);
  assign _zz__24_10_inner_macOut_2 = (($signed(_zz__24_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_10_inner_activation;
    end else begin
      io_macOut = _24_10_inner_macOut;
    end
  end

  assign _zz__24_10_inner_macOut = ($signed(_zz__zz__24_10_inner_macOut) + $signed(_zz__zz__24_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_10_inner_activation <= 8'h00;
      _24_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_10_inner_activation <= io_addInput;
      end else begin
        _24_10_inner_macOut <= _zz__24_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_777 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_9_inner_macOut;
  wire       [15:0]   _zz__zz__24_9_inner_macOut_1;
  wire       [15:0]   _zz__24_9_inner_macOut_1;
  wire       [15:0]   _zz__24_9_inner_macOut_2;
  reg        [7:0]    _24_9_inner_activation;
  reg        [7:0]    _24_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_9_inner_macOut;

  assign _zz__zz__24_9_inner_macOut = ($signed(io_mulInput) * $signed(_24_9_inner_activation));
  assign _zz__zz__24_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_9_inner_macOut)) ? 16'h007f : _zz__24_9_inner_macOut_2);
  assign _zz__24_9_inner_macOut_2 = (($signed(_zz__24_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_9_inner_activation;
    end else begin
      io_macOut = _24_9_inner_macOut;
    end
  end

  assign _zz__24_9_inner_macOut = ($signed(_zz__zz__24_9_inner_macOut) + $signed(_zz__zz__24_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_9_inner_activation <= 8'h00;
      _24_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_9_inner_activation <= io_addInput;
      end else begin
        _24_9_inner_macOut <= _zz__24_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_776 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_8_inner_macOut;
  wire       [15:0]   _zz__zz__24_8_inner_macOut_1;
  wire       [15:0]   _zz__24_8_inner_macOut_1;
  wire       [15:0]   _zz__24_8_inner_macOut_2;
  reg        [7:0]    _24_8_inner_activation;
  reg        [7:0]    _24_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_8_inner_macOut;

  assign _zz__zz__24_8_inner_macOut = ($signed(io_mulInput) * $signed(_24_8_inner_activation));
  assign _zz__zz__24_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_8_inner_macOut)) ? 16'h007f : _zz__24_8_inner_macOut_2);
  assign _zz__24_8_inner_macOut_2 = (($signed(_zz__24_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_8_inner_activation;
    end else begin
      io_macOut = _24_8_inner_macOut;
    end
  end

  assign _zz__24_8_inner_macOut = ($signed(_zz__zz__24_8_inner_macOut) + $signed(_zz__zz__24_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_8_inner_activation <= 8'h00;
      _24_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_8_inner_activation <= io_addInput;
      end else begin
        _24_8_inner_macOut <= _zz__24_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_775 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_7_inner_macOut;
  wire       [15:0]   _zz__zz__24_7_inner_macOut_1;
  wire       [15:0]   _zz__24_7_inner_macOut_1;
  wire       [15:0]   _zz__24_7_inner_macOut_2;
  reg        [7:0]    _24_7_inner_activation;
  reg        [7:0]    _24_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_7_inner_macOut;

  assign _zz__zz__24_7_inner_macOut = ($signed(io_mulInput) * $signed(_24_7_inner_activation));
  assign _zz__zz__24_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_7_inner_macOut)) ? 16'h007f : _zz__24_7_inner_macOut_2);
  assign _zz__24_7_inner_macOut_2 = (($signed(_zz__24_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_7_inner_activation;
    end else begin
      io_macOut = _24_7_inner_macOut;
    end
  end

  assign _zz__24_7_inner_macOut = ($signed(_zz__zz__24_7_inner_macOut) + $signed(_zz__zz__24_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_7_inner_activation <= 8'h00;
      _24_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_7_inner_activation <= io_addInput;
      end else begin
        _24_7_inner_macOut <= _zz__24_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_774 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_6_inner_macOut;
  wire       [15:0]   _zz__zz__24_6_inner_macOut_1;
  wire       [15:0]   _zz__24_6_inner_macOut_1;
  wire       [15:0]   _zz__24_6_inner_macOut_2;
  reg        [7:0]    _24_6_inner_activation;
  reg        [7:0]    _24_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_6_inner_macOut;

  assign _zz__zz__24_6_inner_macOut = ($signed(io_mulInput) * $signed(_24_6_inner_activation));
  assign _zz__zz__24_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_6_inner_macOut)) ? 16'h007f : _zz__24_6_inner_macOut_2);
  assign _zz__24_6_inner_macOut_2 = (($signed(_zz__24_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_6_inner_activation;
    end else begin
      io_macOut = _24_6_inner_macOut;
    end
  end

  assign _zz__24_6_inner_macOut = ($signed(_zz__zz__24_6_inner_macOut) + $signed(_zz__zz__24_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_6_inner_activation <= 8'h00;
      _24_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_6_inner_activation <= io_addInput;
      end else begin
        _24_6_inner_macOut <= _zz__24_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_773 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_5_inner_macOut;
  wire       [15:0]   _zz__zz__24_5_inner_macOut_1;
  wire       [15:0]   _zz__24_5_inner_macOut_1;
  wire       [15:0]   _zz__24_5_inner_macOut_2;
  reg        [7:0]    _24_5_inner_activation;
  reg        [7:0]    _24_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_5_inner_macOut;

  assign _zz__zz__24_5_inner_macOut = ($signed(io_mulInput) * $signed(_24_5_inner_activation));
  assign _zz__zz__24_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_5_inner_macOut)) ? 16'h007f : _zz__24_5_inner_macOut_2);
  assign _zz__24_5_inner_macOut_2 = (($signed(_zz__24_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_5_inner_activation;
    end else begin
      io_macOut = _24_5_inner_macOut;
    end
  end

  assign _zz__24_5_inner_macOut = ($signed(_zz__zz__24_5_inner_macOut) + $signed(_zz__zz__24_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_5_inner_activation <= 8'h00;
      _24_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_5_inner_activation <= io_addInput;
      end else begin
        _24_5_inner_macOut <= _zz__24_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_772 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_4_inner_macOut;
  wire       [15:0]   _zz__zz__24_4_inner_macOut_1;
  wire       [15:0]   _zz__24_4_inner_macOut_1;
  wire       [15:0]   _zz__24_4_inner_macOut_2;
  reg        [7:0]    _24_4_inner_activation;
  reg        [7:0]    _24_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_4_inner_macOut;

  assign _zz__zz__24_4_inner_macOut = ($signed(io_mulInput) * $signed(_24_4_inner_activation));
  assign _zz__zz__24_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_4_inner_macOut)) ? 16'h007f : _zz__24_4_inner_macOut_2);
  assign _zz__24_4_inner_macOut_2 = (($signed(_zz__24_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_4_inner_activation;
    end else begin
      io_macOut = _24_4_inner_macOut;
    end
  end

  assign _zz__24_4_inner_macOut = ($signed(_zz__zz__24_4_inner_macOut) + $signed(_zz__zz__24_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_4_inner_activation <= 8'h00;
      _24_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_4_inner_activation <= io_addInput;
      end else begin
        _24_4_inner_macOut <= _zz__24_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_771 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_3_inner_macOut;
  wire       [15:0]   _zz__zz__24_3_inner_macOut_1;
  wire       [15:0]   _zz__24_3_inner_macOut_1;
  wire       [15:0]   _zz__24_3_inner_macOut_2;
  reg        [7:0]    _24_3_inner_activation;
  reg        [7:0]    _24_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_3_inner_macOut;

  assign _zz__zz__24_3_inner_macOut = ($signed(io_mulInput) * $signed(_24_3_inner_activation));
  assign _zz__zz__24_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_3_inner_macOut)) ? 16'h007f : _zz__24_3_inner_macOut_2);
  assign _zz__24_3_inner_macOut_2 = (($signed(_zz__24_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_3_inner_activation;
    end else begin
      io_macOut = _24_3_inner_macOut;
    end
  end

  assign _zz__24_3_inner_macOut = ($signed(_zz__zz__24_3_inner_macOut) + $signed(_zz__zz__24_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_3_inner_activation <= 8'h00;
      _24_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_3_inner_activation <= io_addInput;
      end else begin
        _24_3_inner_macOut <= _zz__24_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_770 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_2_inner_macOut;
  wire       [15:0]   _zz__zz__24_2_inner_macOut_1;
  wire       [15:0]   _zz__24_2_inner_macOut_1;
  wire       [15:0]   _zz__24_2_inner_macOut_2;
  reg        [7:0]    _24_2_inner_activation;
  reg        [7:0]    _24_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_2_inner_macOut;

  assign _zz__zz__24_2_inner_macOut = ($signed(io_mulInput) * $signed(_24_2_inner_activation));
  assign _zz__zz__24_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_2_inner_macOut)) ? 16'h007f : _zz__24_2_inner_macOut_2);
  assign _zz__24_2_inner_macOut_2 = (($signed(_zz__24_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_2_inner_activation;
    end else begin
      io_macOut = _24_2_inner_macOut;
    end
  end

  assign _zz__24_2_inner_macOut = ($signed(_zz__zz__24_2_inner_macOut) + $signed(_zz__zz__24_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_2_inner_activation <= 8'h00;
      _24_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_2_inner_activation <= io_addInput;
      end else begin
        _24_2_inner_macOut <= _zz__24_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_769 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_1_inner_macOut;
  wire       [15:0]   _zz__zz__24_1_inner_macOut_1;
  wire       [15:0]   _zz__24_1_inner_macOut_1;
  wire       [15:0]   _zz__24_1_inner_macOut_2;
  reg        [7:0]    _24_1_inner_activation;
  reg        [7:0]    _24_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_1_inner_macOut;

  assign _zz__zz__24_1_inner_macOut = ($signed(io_mulInput) * $signed(_24_1_inner_activation));
  assign _zz__zz__24_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_1_inner_macOut)) ? 16'h007f : _zz__24_1_inner_macOut_2);
  assign _zz__24_1_inner_macOut_2 = (($signed(_zz__24_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_1_inner_activation;
    end else begin
      io_macOut = _24_1_inner_macOut;
    end
  end

  assign _zz__24_1_inner_macOut = ($signed(_zz__zz__24_1_inner_macOut) + $signed(_zz__zz__24_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_1_inner_activation <= 8'h00;
      _24_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_1_inner_activation <= io_addInput;
      end else begin
        _24_1_inner_macOut <= _zz__24_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_768 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__24_0_inner_macOut;
  wire       [15:0]   _zz__zz__24_0_inner_macOut_1;
  wire       [15:0]   _zz__24_0_inner_macOut_1;
  wire       [15:0]   _zz__24_0_inner_macOut_2;
  reg        [7:0]    _24_0_inner_activation;
  reg        [7:0]    _24_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__24_0_inner_macOut;

  assign _zz__zz__24_0_inner_macOut = ($signed(io_mulInput) * $signed(_24_0_inner_activation));
  assign _zz__zz__24_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__24_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__24_0_inner_macOut)) ? 16'h007f : _zz__24_0_inner_macOut_2);
  assign _zz__24_0_inner_macOut_2 = (($signed(_zz__24_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__24_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _24_0_inner_activation;
    end else begin
      io_macOut = _24_0_inner_macOut;
    end
  end

  assign _zz__24_0_inner_macOut = ($signed(_zz__zz__24_0_inner_macOut) + $signed(_zz__zz__24_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _24_0_inner_activation <= 8'h00;
      _24_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _24_0_inner_activation <= io_addInput;
      end else begin
        _24_0_inner_macOut <= _zz__24_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_767 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_31_inner_macOut;
  wire       [15:0]   _zz__zz__23_31_inner_macOut_1;
  wire       [15:0]   _zz__23_31_inner_macOut_1;
  wire       [15:0]   _zz__23_31_inner_macOut_2;
  reg        [7:0]    _23_31_inner_activation;
  reg        [7:0]    _23_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_31_inner_macOut;

  assign _zz__zz__23_31_inner_macOut = ($signed(io_mulInput) * $signed(_23_31_inner_activation));
  assign _zz__zz__23_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_31_inner_macOut)) ? 16'h007f : _zz__23_31_inner_macOut_2);
  assign _zz__23_31_inner_macOut_2 = (($signed(_zz__23_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_31_inner_activation;
    end else begin
      io_macOut = _23_31_inner_macOut;
    end
  end

  assign _zz__23_31_inner_macOut = ($signed(_zz__zz__23_31_inner_macOut) + $signed(_zz__zz__23_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_31_inner_activation <= 8'h00;
      _23_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_31_inner_activation <= io_addInput;
      end else begin
        _23_31_inner_macOut <= _zz__23_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_766 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_30_inner_macOut;
  wire       [15:0]   _zz__zz__23_30_inner_macOut_1;
  wire       [15:0]   _zz__23_30_inner_macOut_1;
  wire       [15:0]   _zz__23_30_inner_macOut_2;
  reg        [7:0]    _23_30_inner_activation;
  reg        [7:0]    _23_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_30_inner_macOut;

  assign _zz__zz__23_30_inner_macOut = ($signed(io_mulInput) * $signed(_23_30_inner_activation));
  assign _zz__zz__23_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_30_inner_macOut)) ? 16'h007f : _zz__23_30_inner_macOut_2);
  assign _zz__23_30_inner_macOut_2 = (($signed(_zz__23_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_30_inner_activation;
    end else begin
      io_macOut = _23_30_inner_macOut;
    end
  end

  assign _zz__23_30_inner_macOut = ($signed(_zz__zz__23_30_inner_macOut) + $signed(_zz__zz__23_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_30_inner_activation <= 8'h00;
      _23_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_30_inner_activation <= io_addInput;
      end else begin
        _23_30_inner_macOut <= _zz__23_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_765 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_29_inner_macOut;
  wire       [15:0]   _zz__zz__23_29_inner_macOut_1;
  wire       [15:0]   _zz__23_29_inner_macOut_1;
  wire       [15:0]   _zz__23_29_inner_macOut_2;
  reg        [7:0]    _23_29_inner_activation;
  reg        [7:0]    _23_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_29_inner_macOut;

  assign _zz__zz__23_29_inner_macOut = ($signed(io_mulInput) * $signed(_23_29_inner_activation));
  assign _zz__zz__23_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_29_inner_macOut)) ? 16'h007f : _zz__23_29_inner_macOut_2);
  assign _zz__23_29_inner_macOut_2 = (($signed(_zz__23_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_29_inner_activation;
    end else begin
      io_macOut = _23_29_inner_macOut;
    end
  end

  assign _zz__23_29_inner_macOut = ($signed(_zz__zz__23_29_inner_macOut) + $signed(_zz__zz__23_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_29_inner_activation <= 8'h00;
      _23_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_29_inner_activation <= io_addInput;
      end else begin
        _23_29_inner_macOut <= _zz__23_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_764 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_28_inner_macOut;
  wire       [15:0]   _zz__zz__23_28_inner_macOut_1;
  wire       [15:0]   _zz__23_28_inner_macOut_1;
  wire       [15:0]   _zz__23_28_inner_macOut_2;
  reg        [7:0]    _23_28_inner_activation;
  reg        [7:0]    _23_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_28_inner_macOut;

  assign _zz__zz__23_28_inner_macOut = ($signed(io_mulInput) * $signed(_23_28_inner_activation));
  assign _zz__zz__23_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_28_inner_macOut)) ? 16'h007f : _zz__23_28_inner_macOut_2);
  assign _zz__23_28_inner_macOut_2 = (($signed(_zz__23_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_28_inner_activation;
    end else begin
      io_macOut = _23_28_inner_macOut;
    end
  end

  assign _zz__23_28_inner_macOut = ($signed(_zz__zz__23_28_inner_macOut) + $signed(_zz__zz__23_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_28_inner_activation <= 8'h00;
      _23_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_28_inner_activation <= io_addInput;
      end else begin
        _23_28_inner_macOut <= _zz__23_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_763 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_27_inner_macOut;
  wire       [15:0]   _zz__zz__23_27_inner_macOut_1;
  wire       [15:0]   _zz__23_27_inner_macOut_1;
  wire       [15:0]   _zz__23_27_inner_macOut_2;
  reg        [7:0]    _23_27_inner_activation;
  reg        [7:0]    _23_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_27_inner_macOut;

  assign _zz__zz__23_27_inner_macOut = ($signed(io_mulInput) * $signed(_23_27_inner_activation));
  assign _zz__zz__23_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_27_inner_macOut)) ? 16'h007f : _zz__23_27_inner_macOut_2);
  assign _zz__23_27_inner_macOut_2 = (($signed(_zz__23_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_27_inner_activation;
    end else begin
      io_macOut = _23_27_inner_macOut;
    end
  end

  assign _zz__23_27_inner_macOut = ($signed(_zz__zz__23_27_inner_macOut) + $signed(_zz__zz__23_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_27_inner_activation <= 8'h00;
      _23_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_27_inner_activation <= io_addInput;
      end else begin
        _23_27_inner_macOut <= _zz__23_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_762 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_26_inner_macOut;
  wire       [15:0]   _zz__zz__23_26_inner_macOut_1;
  wire       [15:0]   _zz__23_26_inner_macOut_1;
  wire       [15:0]   _zz__23_26_inner_macOut_2;
  reg        [7:0]    _23_26_inner_activation;
  reg        [7:0]    _23_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_26_inner_macOut;

  assign _zz__zz__23_26_inner_macOut = ($signed(io_mulInput) * $signed(_23_26_inner_activation));
  assign _zz__zz__23_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_26_inner_macOut)) ? 16'h007f : _zz__23_26_inner_macOut_2);
  assign _zz__23_26_inner_macOut_2 = (($signed(_zz__23_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_26_inner_activation;
    end else begin
      io_macOut = _23_26_inner_macOut;
    end
  end

  assign _zz__23_26_inner_macOut = ($signed(_zz__zz__23_26_inner_macOut) + $signed(_zz__zz__23_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_26_inner_activation <= 8'h00;
      _23_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_26_inner_activation <= io_addInput;
      end else begin
        _23_26_inner_macOut <= _zz__23_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_761 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_25_inner_macOut;
  wire       [15:0]   _zz__zz__23_25_inner_macOut_1;
  wire       [15:0]   _zz__23_25_inner_macOut_1;
  wire       [15:0]   _zz__23_25_inner_macOut_2;
  reg        [7:0]    _23_25_inner_activation;
  reg        [7:0]    _23_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_25_inner_macOut;

  assign _zz__zz__23_25_inner_macOut = ($signed(io_mulInput) * $signed(_23_25_inner_activation));
  assign _zz__zz__23_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_25_inner_macOut)) ? 16'h007f : _zz__23_25_inner_macOut_2);
  assign _zz__23_25_inner_macOut_2 = (($signed(_zz__23_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_25_inner_activation;
    end else begin
      io_macOut = _23_25_inner_macOut;
    end
  end

  assign _zz__23_25_inner_macOut = ($signed(_zz__zz__23_25_inner_macOut) + $signed(_zz__zz__23_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_25_inner_activation <= 8'h00;
      _23_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_25_inner_activation <= io_addInput;
      end else begin
        _23_25_inner_macOut <= _zz__23_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_760 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_24_inner_macOut;
  wire       [15:0]   _zz__zz__23_24_inner_macOut_1;
  wire       [15:0]   _zz__23_24_inner_macOut_1;
  wire       [15:0]   _zz__23_24_inner_macOut_2;
  reg        [7:0]    _23_24_inner_activation;
  reg        [7:0]    _23_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_24_inner_macOut;

  assign _zz__zz__23_24_inner_macOut = ($signed(io_mulInput) * $signed(_23_24_inner_activation));
  assign _zz__zz__23_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_24_inner_macOut)) ? 16'h007f : _zz__23_24_inner_macOut_2);
  assign _zz__23_24_inner_macOut_2 = (($signed(_zz__23_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_24_inner_activation;
    end else begin
      io_macOut = _23_24_inner_macOut;
    end
  end

  assign _zz__23_24_inner_macOut = ($signed(_zz__zz__23_24_inner_macOut) + $signed(_zz__zz__23_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_24_inner_activation <= 8'h00;
      _23_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_24_inner_activation <= io_addInput;
      end else begin
        _23_24_inner_macOut <= _zz__23_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_759 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_23_inner_macOut;
  wire       [15:0]   _zz__zz__23_23_inner_macOut_1;
  wire       [15:0]   _zz__23_23_inner_macOut_1;
  wire       [15:0]   _zz__23_23_inner_macOut_2;
  reg        [7:0]    _23_23_inner_activation;
  reg        [7:0]    _23_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_23_inner_macOut;

  assign _zz__zz__23_23_inner_macOut = ($signed(io_mulInput) * $signed(_23_23_inner_activation));
  assign _zz__zz__23_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_23_inner_macOut)) ? 16'h007f : _zz__23_23_inner_macOut_2);
  assign _zz__23_23_inner_macOut_2 = (($signed(_zz__23_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_23_inner_activation;
    end else begin
      io_macOut = _23_23_inner_macOut;
    end
  end

  assign _zz__23_23_inner_macOut = ($signed(_zz__zz__23_23_inner_macOut) + $signed(_zz__zz__23_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_23_inner_activation <= 8'h00;
      _23_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_23_inner_activation <= io_addInput;
      end else begin
        _23_23_inner_macOut <= _zz__23_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_758 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_22_inner_macOut;
  wire       [15:0]   _zz__zz__23_22_inner_macOut_1;
  wire       [15:0]   _zz__23_22_inner_macOut_1;
  wire       [15:0]   _zz__23_22_inner_macOut_2;
  reg        [7:0]    _23_22_inner_activation;
  reg        [7:0]    _23_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_22_inner_macOut;

  assign _zz__zz__23_22_inner_macOut = ($signed(io_mulInput) * $signed(_23_22_inner_activation));
  assign _zz__zz__23_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_22_inner_macOut)) ? 16'h007f : _zz__23_22_inner_macOut_2);
  assign _zz__23_22_inner_macOut_2 = (($signed(_zz__23_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_22_inner_activation;
    end else begin
      io_macOut = _23_22_inner_macOut;
    end
  end

  assign _zz__23_22_inner_macOut = ($signed(_zz__zz__23_22_inner_macOut) + $signed(_zz__zz__23_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_22_inner_activation <= 8'h00;
      _23_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_22_inner_activation <= io_addInput;
      end else begin
        _23_22_inner_macOut <= _zz__23_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_757 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_21_inner_macOut;
  wire       [15:0]   _zz__zz__23_21_inner_macOut_1;
  wire       [15:0]   _zz__23_21_inner_macOut_1;
  wire       [15:0]   _zz__23_21_inner_macOut_2;
  reg        [7:0]    _23_21_inner_activation;
  reg        [7:0]    _23_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_21_inner_macOut;

  assign _zz__zz__23_21_inner_macOut = ($signed(io_mulInput) * $signed(_23_21_inner_activation));
  assign _zz__zz__23_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_21_inner_macOut)) ? 16'h007f : _zz__23_21_inner_macOut_2);
  assign _zz__23_21_inner_macOut_2 = (($signed(_zz__23_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_21_inner_activation;
    end else begin
      io_macOut = _23_21_inner_macOut;
    end
  end

  assign _zz__23_21_inner_macOut = ($signed(_zz__zz__23_21_inner_macOut) + $signed(_zz__zz__23_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_21_inner_activation <= 8'h00;
      _23_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_21_inner_activation <= io_addInput;
      end else begin
        _23_21_inner_macOut <= _zz__23_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_756 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_20_inner_macOut;
  wire       [15:0]   _zz__zz__23_20_inner_macOut_1;
  wire       [15:0]   _zz__23_20_inner_macOut_1;
  wire       [15:0]   _zz__23_20_inner_macOut_2;
  reg        [7:0]    _23_20_inner_activation;
  reg        [7:0]    _23_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_20_inner_macOut;

  assign _zz__zz__23_20_inner_macOut = ($signed(io_mulInput) * $signed(_23_20_inner_activation));
  assign _zz__zz__23_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_20_inner_macOut)) ? 16'h007f : _zz__23_20_inner_macOut_2);
  assign _zz__23_20_inner_macOut_2 = (($signed(_zz__23_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_20_inner_activation;
    end else begin
      io_macOut = _23_20_inner_macOut;
    end
  end

  assign _zz__23_20_inner_macOut = ($signed(_zz__zz__23_20_inner_macOut) + $signed(_zz__zz__23_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_20_inner_activation <= 8'h00;
      _23_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_20_inner_activation <= io_addInput;
      end else begin
        _23_20_inner_macOut <= _zz__23_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_755 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_19_inner_macOut;
  wire       [15:0]   _zz__zz__23_19_inner_macOut_1;
  wire       [15:0]   _zz__23_19_inner_macOut_1;
  wire       [15:0]   _zz__23_19_inner_macOut_2;
  reg        [7:0]    _23_19_inner_activation;
  reg        [7:0]    _23_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_19_inner_macOut;

  assign _zz__zz__23_19_inner_macOut = ($signed(io_mulInput) * $signed(_23_19_inner_activation));
  assign _zz__zz__23_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_19_inner_macOut)) ? 16'h007f : _zz__23_19_inner_macOut_2);
  assign _zz__23_19_inner_macOut_2 = (($signed(_zz__23_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_19_inner_activation;
    end else begin
      io_macOut = _23_19_inner_macOut;
    end
  end

  assign _zz__23_19_inner_macOut = ($signed(_zz__zz__23_19_inner_macOut) + $signed(_zz__zz__23_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_19_inner_activation <= 8'h00;
      _23_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_19_inner_activation <= io_addInput;
      end else begin
        _23_19_inner_macOut <= _zz__23_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_754 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_18_inner_macOut;
  wire       [15:0]   _zz__zz__23_18_inner_macOut_1;
  wire       [15:0]   _zz__23_18_inner_macOut_1;
  wire       [15:0]   _zz__23_18_inner_macOut_2;
  reg        [7:0]    _23_18_inner_activation;
  reg        [7:0]    _23_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_18_inner_macOut;

  assign _zz__zz__23_18_inner_macOut = ($signed(io_mulInput) * $signed(_23_18_inner_activation));
  assign _zz__zz__23_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_18_inner_macOut)) ? 16'h007f : _zz__23_18_inner_macOut_2);
  assign _zz__23_18_inner_macOut_2 = (($signed(_zz__23_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_18_inner_activation;
    end else begin
      io_macOut = _23_18_inner_macOut;
    end
  end

  assign _zz__23_18_inner_macOut = ($signed(_zz__zz__23_18_inner_macOut) + $signed(_zz__zz__23_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_18_inner_activation <= 8'h00;
      _23_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_18_inner_activation <= io_addInput;
      end else begin
        _23_18_inner_macOut <= _zz__23_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_753 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_17_inner_macOut;
  wire       [15:0]   _zz__zz__23_17_inner_macOut_1;
  wire       [15:0]   _zz__23_17_inner_macOut_1;
  wire       [15:0]   _zz__23_17_inner_macOut_2;
  reg        [7:0]    _23_17_inner_activation;
  reg        [7:0]    _23_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_17_inner_macOut;

  assign _zz__zz__23_17_inner_macOut = ($signed(io_mulInput) * $signed(_23_17_inner_activation));
  assign _zz__zz__23_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_17_inner_macOut)) ? 16'h007f : _zz__23_17_inner_macOut_2);
  assign _zz__23_17_inner_macOut_2 = (($signed(_zz__23_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_17_inner_activation;
    end else begin
      io_macOut = _23_17_inner_macOut;
    end
  end

  assign _zz__23_17_inner_macOut = ($signed(_zz__zz__23_17_inner_macOut) + $signed(_zz__zz__23_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_17_inner_activation <= 8'h00;
      _23_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_17_inner_activation <= io_addInput;
      end else begin
        _23_17_inner_macOut <= _zz__23_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_752 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_16_inner_macOut;
  wire       [15:0]   _zz__zz__23_16_inner_macOut_1;
  wire       [15:0]   _zz__23_16_inner_macOut_1;
  wire       [15:0]   _zz__23_16_inner_macOut_2;
  reg        [7:0]    _23_16_inner_activation;
  reg        [7:0]    _23_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_16_inner_macOut;

  assign _zz__zz__23_16_inner_macOut = ($signed(io_mulInput) * $signed(_23_16_inner_activation));
  assign _zz__zz__23_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_16_inner_macOut)) ? 16'h007f : _zz__23_16_inner_macOut_2);
  assign _zz__23_16_inner_macOut_2 = (($signed(_zz__23_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_16_inner_activation;
    end else begin
      io_macOut = _23_16_inner_macOut;
    end
  end

  assign _zz__23_16_inner_macOut = ($signed(_zz__zz__23_16_inner_macOut) + $signed(_zz__zz__23_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_16_inner_activation <= 8'h00;
      _23_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_16_inner_activation <= io_addInput;
      end else begin
        _23_16_inner_macOut <= _zz__23_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_751 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_15_inner_macOut;
  wire       [15:0]   _zz__zz__23_15_inner_macOut_1;
  wire       [15:0]   _zz__23_15_inner_macOut_1;
  wire       [15:0]   _zz__23_15_inner_macOut_2;
  reg        [7:0]    _23_15_inner_activation;
  reg        [7:0]    _23_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_15_inner_macOut;

  assign _zz__zz__23_15_inner_macOut = ($signed(io_mulInput) * $signed(_23_15_inner_activation));
  assign _zz__zz__23_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_15_inner_macOut)) ? 16'h007f : _zz__23_15_inner_macOut_2);
  assign _zz__23_15_inner_macOut_2 = (($signed(_zz__23_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_15_inner_activation;
    end else begin
      io_macOut = _23_15_inner_macOut;
    end
  end

  assign _zz__23_15_inner_macOut = ($signed(_zz__zz__23_15_inner_macOut) + $signed(_zz__zz__23_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_15_inner_activation <= 8'h00;
      _23_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_15_inner_activation <= io_addInput;
      end else begin
        _23_15_inner_macOut <= _zz__23_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_750 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_14_inner_macOut;
  wire       [15:0]   _zz__zz__23_14_inner_macOut_1;
  wire       [15:0]   _zz__23_14_inner_macOut_1;
  wire       [15:0]   _zz__23_14_inner_macOut_2;
  reg        [7:0]    _23_14_inner_activation;
  reg        [7:0]    _23_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_14_inner_macOut;

  assign _zz__zz__23_14_inner_macOut = ($signed(io_mulInput) * $signed(_23_14_inner_activation));
  assign _zz__zz__23_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_14_inner_macOut)) ? 16'h007f : _zz__23_14_inner_macOut_2);
  assign _zz__23_14_inner_macOut_2 = (($signed(_zz__23_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_14_inner_activation;
    end else begin
      io_macOut = _23_14_inner_macOut;
    end
  end

  assign _zz__23_14_inner_macOut = ($signed(_zz__zz__23_14_inner_macOut) + $signed(_zz__zz__23_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_14_inner_activation <= 8'h00;
      _23_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_14_inner_activation <= io_addInput;
      end else begin
        _23_14_inner_macOut <= _zz__23_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_749 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_13_inner_macOut;
  wire       [15:0]   _zz__zz__23_13_inner_macOut_1;
  wire       [15:0]   _zz__23_13_inner_macOut_1;
  wire       [15:0]   _zz__23_13_inner_macOut_2;
  reg        [7:0]    _23_13_inner_activation;
  reg        [7:0]    _23_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_13_inner_macOut;

  assign _zz__zz__23_13_inner_macOut = ($signed(io_mulInput) * $signed(_23_13_inner_activation));
  assign _zz__zz__23_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_13_inner_macOut)) ? 16'h007f : _zz__23_13_inner_macOut_2);
  assign _zz__23_13_inner_macOut_2 = (($signed(_zz__23_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_13_inner_activation;
    end else begin
      io_macOut = _23_13_inner_macOut;
    end
  end

  assign _zz__23_13_inner_macOut = ($signed(_zz__zz__23_13_inner_macOut) + $signed(_zz__zz__23_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_13_inner_activation <= 8'h00;
      _23_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_13_inner_activation <= io_addInput;
      end else begin
        _23_13_inner_macOut <= _zz__23_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_748 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_12_inner_macOut;
  wire       [15:0]   _zz__zz__23_12_inner_macOut_1;
  wire       [15:0]   _zz__23_12_inner_macOut_1;
  wire       [15:0]   _zz__23_12_inner_macOut_2;
  reg        [7:0]    _23_12_inner_activation;
  reg        [7:0]    _23_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_12_inner_macOut;

  assign _zz__zz__23_12_inner_macOut = ($signed(io_mulInput) * $signed(_23_12_inner_activation));
  assign _zz__zz__23_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_12_inner_macOut)) ? 16'h007f : _zz__23_12_inner_macOut_2);
  assign _zz__23_12_inner_macOut_2 = (($signed(_zz__23_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_12_inner_activation;
    end else begin
      io_macOut = _23_12_inner_macOut;
    end
  end

  assign _zz__23_12_inner_macOut = ($signed(_zz__zz__23_12_inner_macOut) + $signed(_zz__zz__23_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_12_inner_activation <= 8'h00;
      _23_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_12_inner_activation <= io_addInput;
      end else begin
        _23_12_inner_macOut <= _zz__23_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_747 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_11_inner_macOut;
  wire       [15:0]   _zz__zz__23_11_inner_macOut_1;
  wire       [15:0]   _zz__23_11_inner_macOut_1;
  wire       [15:0]   _zz__23_11_inner_macOut_2;
  reg        [7:0]    _23_11_inner_activation;
  reg        [7:0]    _23_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_11_inner_macOut;

  assign _zz__zz__23_11_inner_macOut = ($signed(io_mulInput) * $signed(_23_11_inner_activation));
  assign _zz__zz__23_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_11_inner_macOut)) ? 16'h007f : _zz__23_11_inner_macOut_2);
  assign _zz__23_11_inner_macOut_2 = (($signed(_zz__23_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_11_inner_activation;
    end else begin
      io_macOut = _23_11_inner_macOut;
    end
  end

  assign _zz__23_11_inner_macOut = ($signed(_zz__zz__23_11_inner_macOut) + $signed(_zz__zz__23_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_11_inner_activation <= 8'h00;
      _23_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_11_inner_activation <= io_addInput;
      end else begin
        _23_11_inner_macOut <= _zz__23_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_746 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_10_inner_macOut;
  wire       [15:0]   _zz__zz__23_10_inner_macOut_1;
  wire       [15:0]   _zz__23_10_inner_macOut_1;
  wire       [15:0]   _zz__23_10_inner_macOut_2;
  reg        [7:0]    _23_10_inner_activation;
  reg        [7:0]    _23_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_10_inner_macOut;

  assign _zz__zz__23_10_inner_macOut = ($signed(io_mulInput) * $signed(_23_10_inner_activation));
  assign _zz__zz__23_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_10_inner_macOut)) ? 16'h007f : _zz__23_10_inner_macOut_2);
  assign _zz__23_10_inner_macOut_2 = (($signed(_zz__23_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_10_inner_activation;
    end else begin
      io_macOut = _23_10_inner_macOut;
    end
  end

  assign _zz__23_10_inner_macOut = ($signed(_zz__zz__23_10_inner_macOut) + $signed(_zz__zz__23_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_10_inner_activation <= 8'h00;
      _23_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_10_inner_activation <= io_addInput;
      end else begin
        _23_10_inner_macOut <= _zz__23_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_745 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_9_inner_macOut;
  wire       [15:0]   _zz__zz__23_9_inner_macOut_1;
  wire       [15:0]   _zz__23_9_inner_macOut_1;
  wire       [15:0]   _zz__23_9_inner_macOut_2;
  reg        [7:0]    _23_9_inner_activation;
  reg        [7:0]    _23_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_9_inner_macOut;

  assign _zz__zz__23_9_inner_macOut = ($signed(io_mulInput) * $signed(_23_9_inner_activation));
  assign _zz__zz__23_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_9_inner_macOut)) ? 16'h007f : _zz__23_9_inner_macOut_2);
  assign _zz__23_9_inner_macOut_2 = (($signed(_zz__23_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_9_inner_activation;
    end else begin
      io_macOut = _23_9_inner_macOut;
    end
  end

  assign _zz__23_9_inner_macOut = ($signed(_zz__zz__23_9_inner_macOut) + $signed(_zz__zz__23_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_9_inner_activation <= 8'h00;
      _23_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_9_inner_activation <= io_addInput;
      end else begin
        _23_9_inner_macOut <= _zz__23_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_744 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_8_inner_macOut;
  wire       [15:0]   _zz__zz__23_8_inner_macOut_1;
  wire       [15:0]   _zz__23_8_inner_macOut_1;
  wire       [15:0]   _zz__23_8_inner_macOut_2;
  reg        [7:0]    _23_8_inner_activation;
  reg        [7:0]    _23_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_8_inner_macOut;

  assign _zz__zz__23_8_inner_macOut = ($signed(io_mulInput) * $signed(_23_8_inner_activation));
  assign _zz__zz__23_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_8_inner_macOut)) ? 16'h007f : _zz__23_8_inner_macOut_2);
  assign _zz__23_8_inner_macOut_2 = (($signed(_zz__23_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_8_inner_activation;
    end else begin
      io_macOut = _23_8_inner_macOut;
    end
  end

  assign _zz__23_8_inner_macOut = ($signed(_zz__zz__23_8_inner_macOut) + $signed(_zz__zz__23_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_8_inner_activation <= 8'h00;
      _23_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_8_inner_activation <= io_addInput;
      end else begin
        _23_8_inner_macOut <= _zz__23_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_743 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_7_inner_macOut;
  wire       [15:0]   _zz__zz__23_7_inner_macOut_1;
  wire       [15:0]   _zz__23_7_inner_macOut_1;
  wire       [15:0]   _zz__23_7_inner_macOut_2;
  reg        [7:0]    _23_7_inner_activation;
  reg        [7:0]    _23_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_7_inner_macOut;

  assign _zz__zz__23_7_inner_macOut = ($signed(io_mulInput) * $signed(_23_7_inner_activation));
  assign _zz__zz__23_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_7_inner_macOut)) ? 16'h007f : _zz__23_7_inner_macOut_2);
  assign _zz__23_7_inner_macOut_2 = (($signed(_zz__23_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_7_inner_activation;
    end else begin
      io_macOut = _23_7_inner_macOut;
    end
  end

  assign _zz__23_7_inner_macOut = ($signed(_zz__zz__23_7_inner_macOut) + $signed(_zz__zz__23_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_7_inner_activation <= 8'h00;
      _23_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_7_inner_activation <= io_addInput;
      end else begin
        _23_7_inner_macOut <= _zz__23_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_742 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_6_inner_macOut;
  wire       [15:0]   _zz__zz__23_6_inner_macOut_1;
  wire       [15:0]   _zz__23_6_inner_macOut_1;
  wire       [15:0]   _zz__23_6_inner_macOut_2;
  reg        [7:0]    _23_6_inner_activation;
  reg        [7:0]    _23_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_6_inner_macOut;

  assign _zz__zz__23_6_inner_macOut = ($signed(io_mulInput) * $signed(_23_6_inner_activation));
  assign _zz__zz__23_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_6_inner_macOut)) ? 16'h007f : _zz__23_6_inner_macOut_2);
  assign _zz__23_6_inner_macOut_2 = (($signed(_zz__23_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_6_inner_activation;
    end else begin
      io_macOut = _23_6_inner_macOut;
    end
  end

  assign _zz__23_6_inner_macOut = ($signed(_zz__zz__23_6_inner_macOut) + $signed(_zz__zz__23_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_6_inner_activation <= 8'h00;
      _23_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_6_inner_activation <= io_addInput;
      end else begin
        _23_6_inner_macOut <= _zz__23_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_741 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_5_inner_macOut;
  wire       [15:0]   _zz__zz__23_5_inner_macOut_1;
  wire       [15:0]   _zz__23_5_inner_macOut_1;
  wire       [15:0]   _zz__23_5_inner_macOut_2;
  reg        [7:0]    _23_5_inner_activation;
  reg        [7:0]    _23_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_5_inner_macOut;

  assign _zz__zz__23_5_inner_macOut = ($signed(io_mulInput) * $signed(_23_5_inner_activation));
  assign _zz__zz__23_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_5_inner_macOut)) ? 16'h007f : _zz__23_5_inner_macOut_2);
  assign _zz__23_5_inner_macOut_2 = (($signed(_zz__23_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_5_inner_activation;
    end else begin
      io_macOut = _23_5_inner_macOut;
    end
  end

  assign _zz__23_5_inner_macOut = ($signed(_zz__zz__23_5_inner_macOut) + $signed(_zz__zz__23_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_5_inner_activation <= 8'h00;
      _23_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_5_inner_activation <= io_addInput;
      end else begin
        _23_5_inner_macOut <= _zz__23_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_740 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_4_inner_macOut;
  wire       [15:0]   _zz__zz__23_4_inner_macOut_1;
  wire       [15:0]   _zz__23_4_inner_macOut_1;
  wire       [15:0]   _zz__23_4_inner_macOut_2;
  reg        [7:0]    _23_4_inner_activation;
  reg        [7:0]    _23_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_4_inner_macOut;

  assign _zz__zz__23_4_inner_macOut = ($signed(io_mulInput) * $signed(_23_4_inner_activation));
  assign _zz__zz__23_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_4_inner_macOut)) ? 16'h007f : _zz__23_4_inner_macOut_2);
  assign _zz__23_4_inner_macOut_2 = (($signed(_zz__23_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_4_inner_activation;
    end else begin
      io_macOut = _23_4_inner_macOut;
    end
  end

  assign _zz__23_4_inner_macOut = ($signed(_zz__zz__23_4_inner_macOut) + $signed(_zz__zz__23_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_4_inner_activation <= 8'h00;
      _23_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_4_inner_activation <= io_addInput;
      end else begin
        _23_4_inner_macOut <= _zz__23_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_739 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_3_inner_macOut;
  wire       [15:0]   _zz__zz__23_3_inner_macOut_1;
  wire       [15:0]   _zz__23_3_inner_macOut_1;
  wire       [15:0]   _zz__23_3_inner_macOut_2;
  reg        [7:0]    _23_3_inner_activation;
  reg        [7:0]    _23_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_3_inner_macOut;

  assign _zz__zz__23_3_inner_macOut = ($signed(io_mulInput) * $signed(_23_3_inner_activation));
  assign _zz__zz__23_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_3_inner_macOut)) ? 16'h007f : _zz__23_3_inner_macOut_2);
  assign _zz__23_3_inner_macOut_2 = (($signed(_zz__23_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_3_inner_activation;
    end else begin
      io_macOut = _23_3_inner_macOut;
    end
  end

  assign _zz__23_3_inner_macOut = ($signed(_zz__zz__23_3_inner_macOut) + $signed(_zz__zz__23_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_3_inner_activation <= 8'h00;
      _23_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_3_inner_activation <= io_addInput;
      end else begin
        _23_3_inner_macOut <= _zz__23_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_738 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_2_inner_macOut;
  wire       [15:0]   _zz__zz__23_2_inner_macOut_1;
  wire       [15:0]   _zz__23_2_inner_macOut_1;
  wire       [15:0]   _zz__23_2_inner_macOut_2;
  reg        [7:0]    _23_2_inner_activation;
  reg        [7:0]    _23_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_2_inner_macOut;

  assign _zz__zz__23_2_inner_macOut = ($signed(io_mulInput) * $signed(_23_2_inner_activation));
  assign _zz__zz__23_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_2_inner_macOut)) ? 16'h007f : _zz__23_2_inner_macOut_2);
  assign _zz__23_2_inner_macOut_2 = (($signed(_zz__23_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_2_inner_activation;
    end else begin
      io_macOut = _23_2_inner_macOut;
    end
  end

  assign _zz__23_2_inner_macOut = ($signed(_zz__zz__23_2_inner_macOut) + $signed(_zz__zz__23_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_2_inner_activation <= 8'h00;
      _23_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_2_inner_activation <= io_addInput;
      end else begin
        _23_2_inner_macOut <= _zz__23_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_737 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_1_inner_macOut;
  wire       [15:0]   _zz__zz__23_1_inner_macOut_1;
  wire       [15:0]   _zz__23_1_inner_macOut_1;
  wire       [15:0]   _zz__23_1_inner_macOut_2;
  reg        [7:0]    _23_1_inner_activation;
  reg        [7:0]    _23_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_1_inner_macOut;

  assign _zz__zz__23_1_inner_macOut = ($signed(io_mulInput) * $signed(_23_1_inner_activation));
  assign _zz__zz__23_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_1_inner_macOut)) ? 16'h007f : _zz__23_1_inner_macOut_2);
  assign _zz__23_1_inner_macOut_2 = (($signed(_zz__23_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_1_inner_activation;
    end else begin
      io_macOut = _23_1_inner_macOut;
    end
  end

  assign _zz__23_1_inner_macOut = ($signed(_zz__zz__23_1_inner_macOut) + $signed(_zz__zz__23_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_1_inner_activation <= 8'h00;
      _23_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_1_inner_activation <= io_addInput;
      end else begin
        _23_1_inner_macOut <= _zz__23_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_736 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__23_0_inner_macOut;
  wire       [15:0]   _zz__zz__23_0_inner_macOut_1;
  wire       [15:0]   _zz__23_0_inner_macOut_1;
  wire       [15:0]   _zz__23_0_inner_macOut_2;
  reg        [7:0]    _23_0_inner_activation;
  reg        [7:0]    _23_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__23_0_inner_macOut;

  assign _zz__zz__23_0_inner_macOut = ($signed(io_mulInput) * $signed(_23_0_inner_activation));
  assign _zz__zz__23_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__23_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__23_0_inner_macOut)) ? 16'h007f : _zz__23_0_inner_macOut_2);
  assign _zz__23_0_inner_macOut_2 = (($signed(_zz__23_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__23_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _23_0_inner_activation;
    end else begin
      io_macOut = _23_0_inner_macOut;
    end
  end

  assign _zz__23_0_inner_macOut = ($signed(_zz__zz__23_0_inner_macOut) + $signed(_zz__zz__23_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _23_0_inner_activation <= 8'h00;
      _23_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _23_0_inner_activation <= io_addInput;
      end else begin
        _23_0_inner_macOut <= _zz__23_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_735 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_31_inner_macOut;
  wire       [15:0]   _zz__zz__22_31_inner_macOut_1;
  wire       [15:0]   _zz__22_31_inner_macOut_1;
  wire       [15:0]   _zz__22_31_inner_macOut_2;
  reg        [7:0]    _22_31_inner_activation;
  reg        [7:0]    _22_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_31_inner_macOut;

  assign _zz__zz__22_31_inner_macOut = ($signed(io_mulInput) * $signed(_22_31_inner_activation));
  assign _zz__zz__22_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_31_inner_macOut)) ? 16'h007f : _zz__22_31_inner_macOut_2);
  assign _zz__22_31_inner_macOut_2 = (($signed(_zz__22_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_31_inner_activation;
    end else begin
      io_macOut = _22_31_inner_macOut;
    end
  end

  assign _zz__22_31_inner_macOut = ($signed(_zz__zz__22_31_inner_macOut) + $signed(_zz__zz__22_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_31_inner_activation <= 8'h00;
      _22_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_31_inner_activation <= io_addInput;
      end else begin
        _22_31_inner_macOut <= _zz__22_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_734 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_30_inner_macOut;
  wire       [15:0]   _zz__zz__22_30_inner_macOut_1;
  wire       [15:0]   _zz__22_30_inner_macOut_1;
  wire       [15:0]   _zz__22_30_inner_macOut_2;
  reg        [7:0]    _22_30_inner_activation;
  reg        [7:0]    _22_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_30_inner_macOut;

  assign _zz__zz__22_30_inner_macOut = ($signed(io_mulInput) * $signed(_22_30_inner_activation));
  assign _zz__zz__22_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_30_inner_macOut)) ? 16'h007f : _zz__22_30_inner_macOut_2);
  assign _zz__22_30_inner_macOut_2 = (($signed(_zz__22_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_30_inner_activation;
    end else begin
      io_macOut = _22_30_inner_macOut;
    end
  end

  assign _zz__22_30_inner_macOut = ($signed(_zz__zz__22_30_inner_macOut) + $signed(_zz__zz__22_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_30_inner_activation <= 8'h00;
      _22_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_30_inner_activation <= io_addInput;
      end else begin
        _22_30_inner_macOut <= _zz__22_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_733 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_29_inner_macOut;
  wire       [15:0]   _zz__zz__22_29_inner_macOut_1;
  wire       [15:0]   _zz__22_29_inner_macOut_1;
  wire       [15:0]   _zz__22_29_inner_macOut_2;
  reg        [7:0]    _22_29_inner_activation;
  reg        [7:0]    _22_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_29_inner_macOut;

  assign _zz__zz__22_29_inner_macOut = ($signed(io_mulInput) * $signed(_22_29_inner_activation));
  assign _zz__zz__22_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_29_inner_macOut)) ? 16'h007f : _zz__22_29_inner_macOut_2);
  assign _zz__22_29_inner_macOut_2 = (($signed(_zz__22_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_29_inner_activation;
    end else begin
      io_macOut = _22_29_inner_macOut;
    end
  end

  assign _zz__22_29_inner_macOut = ($signed(_zz__zz__22_29_inner_macOut) + $signed(_zz__zz__22_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_29_inner_activation <= 8'h00;
      _22_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_29_inner_activation <= io_addInput;
      end else begin
        _22_29_inner_macOut <= _zz__22_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_732 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_28_inner_macOut;
  wire       [15:0]   _zz__zz__22_28_inner_macOut_1;
  wire       [15:0]   _zz__22_28_inner_macOut_1;
  wire       [15:0]   _zz__22_28_inner_macOut_2;
  reg        [7:0]    _22_28_inner_activation;
  reg        [7:0]    _22_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_28_inner_macOut;

  assign _zz__zz__22_28_inner_macOut = ($signed(io_mulInput) * $signed(_22_28_inner_activation));
  assign _zz__zz__22_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_28_inner_macOut)) ? 16'h007f : _zz__22_28_inner_macOut_2);
  assign _zz__22_28_inner_macOut_2 = (($signed(_zz__22_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_28_inner_activation;
    end else begin
      io_macOut = _22_28_inner_macOut;
    end
  end

  assign _zz__22_28_inner_macOut = ($signed(_zz__zz__22_28_inner_macOut) + $signed(_zz__zz__22_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_28_inner_activation <= 8'h00;
      _22_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_28_inner_activation <= io_addInput;
      end else begin
        _22_28_inner_macOut <= _zz__22_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_731 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_27_inner_macOut;
  wire       [15:0]   _zz__zz__22_27_inner_macOut_1;
  wire       [15:0]   _zz__22_27_inner_macOut_1;
  wire       [15:0]   _zz__22_27_inner_macOut_2;
  reg        [7:0]    _22_27_inner_activation;
  reg        [7:0]    _22_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_27_inner_macOut;

  assign _zz__zz__22_27_inner_macOut = ($signed(io_mulInput) * $signed(_22_27_inner_activation));
  assign _zz__zz__22_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_27_inner_macOut)) ? 16'h007f : _zz__22_27_inner_macOut_2);
  assign _zz__22_27_inner_macOut_2 = (($signed(_zz__22_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_27_inner_activation;
    end else begin
      io_macOut = _22_27_inner_macOut;
    end
  end

  assign _zz__22_27_inner_macOut = ($signed(_zz__zz__22_27_inner_macOut) + $signed(_zz__zz__22_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_27_inner_activation <= 8'h00;
      _22_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_27_inner_activation <= io_addInput;
      end else begin
        _22_27_inner_macOut <= _zz__22_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_730 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_26_inner_macOut;
  wire       [15:0]   _zz__zz__22_26_inner_macOut_1;
  wire       [15:0]   _zz__22_26_inner_macOut_1;
  wire       [15:0]   _zz__22_26_inner_macOut_2;
  reg        [7:0]    _22_26_inner_activation;
  reg        [7:0]    _22_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_26_inner_macOut;

  assign _zz__zz__22_26_inner_macOut = ($signed(io_mulInput) * $signed(_22_26_inner_activation));
  assign _zz__zz__22_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_26_inner_macOut)) ? 16'h007f : _zz__22_26_inner_macOut_2);
  assign _zz__22_26_inner_macOut_2 = (($signed(_zz__22_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_26_inner_activation;
    end else begin
      io_macOut = _22_26_inner_macOut;
    end
  end

  assign _zz__22_26_inner_macOut = ($signed(_zz__zz__22_26_inner_macOut) + $signed(_zz__zz__22_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_26_inner_activation <= 8'h00;
      _22_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_26_inner_activation <= io_addInput;
      end else begin
        _22_26_inner_macOut <= _zz__22_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_729 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_25_inner_macOut;
  wire       [15:0]   _zz__zz__22_25_inner_macOut_1;
  wire       [15:0]   _zz__22_25_inner_macOut_1;
  wire       [15:0]   _zz__22_25_inner_macOut_2;
  reg        [7:0]    _22_25_inner_activation;
  reg        [7:0]    _22_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_25_inner_macOut;

  assign _zz__zz__22_25_inner_macOut = ($signed(io_mulInput) * $signed(_22_25_inner_activation));
  assign _zz__zz__22_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_25_inner_macOut)) ? 16'h007f : _zz__22_25_inner_macOut_2);
  assign _zz__22_25_inner_macOut_2 = (($signed(_zz__22_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_25_inner_activation;
    end else begin
      io_macOut = _22_25_inner_macOut;
    end
  end

  assign _zz__22_25_inner_macOut = ($signed(_zz__zz__22_25_inner_macOut) + $signed(_zz__zz__22_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_25_inner_activation <= 8'h00;
      _22_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_25_inner_activation <= io_addInput;
      end else begin
        _22_25_inner_macOut <= _zz__22_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_728 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_24_inner_macOut;
  wire       [15:0]   _zz__zz__22_24_inner_macOut_1;
  wire       [15:0]   _zz__22_24_inner_macOut_1;
  wire       [15:0]   _zz__22_24_inner_macOut_2;
  reg        [7:0]    _22_24_inner_activation;
  reg        [7:0]    _22_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_24_inner_macOut;

  assign _zz__zz__22_24_inner_macOut = ($signed(io_mulInput) * $signed(_22_24_inner_activation));
  assign _zz__zz__22_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_24_inner_macOut)) ? 16'h007f : _zz__22_24_inner_macOut_2);
  assign _zz__22_24_inner_macOut_2 = (($signed(_zz__22_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_24_inner_activation;
    end else begin
      io_macOut = _22_24_inner_macOut;
    end
  end

  assign _zz__22_24_inner_macOut = ($signed(_zz__zz__22_24_inner_macOut) + $signed(_zz__zz__22_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_24_inner_activation <= 8'h00;
      _22_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_24_inner_activation <= io_addInput;
      end else begin
        _22_24_inner_macOut <= _zz__22_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_727 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_23_inner_macOut;
  wire       [15:0]   _zz__zz__22_23_inner_macOut_1;
  wire       [15:0]   _zz__22_23_inner_macOut_1;
  wire       [15:0]   _zz__22_23_inner_macOut_2;
  reg        [7:0]    _22_23_inner_activation;
  reg        [7:0]    _22_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_23_inner_macOut;

  assign _zz__zz__22_23_inner_macOut = ($signed(io_mulInput) * $signed(_22_23_inner_activation));
  assign _zz__zz__22_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_23_inner_macOut)) ? 16'h007f : _zz__22_23_inner_macOut_2);
  assign _zz__22_23_inner_macOut_2 = (($signed(_zz__22_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_23_inner_activation;
    end else begin
      io_macOut = _22_23_inner_macOut;
    end
  end

  assign _zz__22_23_inner_macOut = ($signed(_zz__zz__22_23_inner_macOut) + $signed(_zz__zz__22_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_23_inner_activation <= 8'h00;
      _22_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_23_inner_activation <= io_addInput;
      end else begin
        _22_23_inner_macOut <= _zz__22_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_726 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_22_inner_macOut;
  wire       [15:0]   _zz__zz__22_22_inner_macOut_1;
  wire       [15:0]   _zz__22_22_inner_macOut_1;
  wire       [15:0]   _zz__22_22_inner_macOut_2;
  reg        [7:0]    _22_22_inner_activation;
  reg        [7:0]    _22_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_22_inner_macOut;

  assign _zz__zz__22_22_inner_macOut = ($signed(io_mulInput) * $signed(_22_22_inner_activation));
  assign _zz__zz__22_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_22_inner_macOut)) ? 16'h007f : _zz__22_22_inner_macOut_2);
  assign _zz__22_22_inner_macOut_2 = (($signed(_zz__22_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_22_inner_activation;
    end else begin
      io_macOut = _22_22_inner_macOut;
    end
  end

  assign _zz__22_22_inner_macOut = ($signed(_zz__zz__22_22_inner_macOut) + $signed(_zz__zz__22_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_22_inner_activation <= 8'h00;
      _22_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_22_inner_activation <= io_addInput;
      end else begin
        _22_22_inner_macOut <= _zz__22_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_725 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_21_inner_macOut;
  wire       [15:0]   _zz__zz__22_21_inner_macOut_1;
  wire       [15:0]   _zz__22_21_inner_macOut_1;
  wire       [15:0]   _zz__22_21_inner_macOut_2;
  reg        [7:0]    _22_21_inner_activation;
  reg        [7:0]    _22_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_21_inner_macOut;

  assign _zz__zz__22_21_inner_macOut = ($signed(io_mulInput) * $signed(_22_21_inner_activation));
  assign _zz__zz__22_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_21_inner_macOut)) ? 16'h007f : _zz__22_21_inner_macOut_2);
  assign _zz__22_21_inner_macOut_2 = (($signed(_zz__22_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_21_inner_activation;
    end else begin
      io_macOut = _22_21_inner_macOut;
    end
  end

  assign _zz__22_21_inner_macOut = ($signed(_zz__zz__22_21_inner_macOut) + $signed(_zz__zz__22_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_21_inner_activation <= 8'h00;
      _22_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_21_inner_activation <= io_addInput;
      end else begin
        _22_21_inner_macOut <= _zz__22_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_724 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_20_inner_macOut;
  wire       [15:0]   _zz__zz__22_20_inner_macOut_1;
  wire       [15:0]   _zz__22_20_inner_macOut_1;
  wire       [15:0]   _zz__22_20_inner_macOut_2;
  reg        [7:0]    _22_20_inner_activation;
  reg        [7:0]    _22_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_20_inner_macOut;

  assign _zz__zz__22_20_inner_macOut = ($signed(io_mulInput) * $signed(_22_20_inner_activation));
  assign _zz__zz__22_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_20_inner_macOut)) ? 16'h007f : _zz__22_20_inner_macOut_2);
  assign _zz__22_20_inner_macOut_2 = (($signed(_zz__22_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_20_inner_activation;
    end else begin
      io_macOut = _22_20_inner_macOut;
    end
  end

  assign _zz__22_20_inner_macOut = ($signed(_zz__zz__22_20_inner_macOut) + $signed(_zz__zz__22_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_20_inner_activation <= 8'h00;
      _22_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_20_inner_activation <= io_addInput;
      end else begin
        _22_20_inner_macOut <= _zz__22_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_723 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_19_inner_macOut;
  wire       [15:0]   _zz__zz__22_19_inner_macOut_1;
  wire       [15:0]   _zz__22_19_inner_macOut_1;
  wire       [15:0]   _zz__22_19_inner_macOut_2;
  reg        [7:0]    _22_19_inner_activation;
  reg        [7:0]    _22_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_19_inner_macOut;

  assign _zz__zz__22_19_inner_macOut = ($signed(io_mulInput) * $signed(_22_19_inner_activation));
  assign _zz__zz__22_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_19_inner_macOut)) ? 16'h007f : _zz__22_19_inner_macOut_2);
  assign _zz__22_19_inner_macOut_2 = (($signed(_zz__22_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_19_inner_activation;
    end else begin
      io_macOut = _22_19_inner_macOut;
    end
  end

  assign _zz__22_19_inner_macOut = ($signed(_zz__zz__22_19_inner_macOut) + $signed(_zz__zz__22_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_19_inner_activation <= 8'h00;
      _22_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_19_inner_activation <= io_addInput;
      end else begin
        _22_19_inner_macOut <= _zz__22_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_722 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_18_inner_macOut;
  wire       [15:0]   _zz__zz__22_18_inner_macOut_1;
  wire       [15:0]   _zz__22_18_inner_macOut_1;
  wire       [15:0]   _zz__22_18_inner_macOut_2;
  reg        [7:0]    _22_18_inner_activation;
  reg        [7:0]    _22_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_18_inner_macOut;

  assign _zz__zz__22_18_inner_macOut = ($signed(io_mulInput) * $signed(_22_18_inner_activation));
  assign _zz__zz__22_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_18_inner_macOut)) ? 16'h007f : _zz__22_18_inner_macOut_2);
  assign _zz__22_18_inner_macOut_2 = (($signed(_zz__22_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_18_inner_activation;
    end else begin
      io_macOut = _22_18_inner_macOut;
    end
  end

  assign _zz__22_18_inner_macOut = ($signed(_zz__zz__22_18_inner_macOut) + $signed(_zz__zz__22_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_18_inner_activation <= 8'h00;
      _22_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_18_inner_activation <= io_addInput;
      end else begin
        _22_18_inner_macOut <= _zz__22_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_721 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_17_inner_macOut;
  wire       [15:0]   _zz__zz__22_17_inner_macOut_1;
  wire       [15:0]   _zz__22_17_inner_macOut_1;
  wire       [15:0]   _zz__22_17_inner_macOut_2;
  reg        [7:0]    _22_17_inner_activation;
  reg        [7:0]    _22_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_17_inner_macOut;

  assign _zz__zz__22_17_inner_macOut = ($signed(io_mulInput) * $signed(_22_17_inner_activation));
  assign _zz__zz__22_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_17_inner_macOut)) ? 16'h007f : _zz__22_17_inner_macOut_2);
  assign _zz__22_17_inner_macOut_2 = (($signed(_zz__22_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_17_inner_activation;
    end else begin
      io_macOut = _22_17_inner_macOut;
    end
  end

  assign _zz__22_17_inner_macOut = ($signed(_zz__zz__22_17_inner_macOut) + $signed(_zz__zz__22_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_17_inner_activation <= 8'h00;
      _22_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_17_inner_activation <= io_addInput;
      end else begin
        _22_17_inner_macOut <= _zz__22_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_720 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_16_inner_macOut;
  wire       [15:0]   _zz__zz__22_16_inner_macOut_1;
  wire       [15:0]   _zz__22_16_inner_macOut_1;
  wire       [15:0]   _zz__22_16_inner_macOut_2;
  reg        [7:0]    _22_16_inner_activation;
  reg        [7:0]    _22_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_16_inner_macOut;

  assign _zz__zz__22_16_inner_macOut = ($signed(io_mulInput) * $signed(_22_16_inner_activation));
  assign _zz__zz__22_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_16_inner_macOut)) ? 16'h007f : _zz__22_16_inner_macOut_2);
  assign _zz__22_16_inner_macOut_2 = (($signed(_zz__22_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_16_inner_activation;
    end else begin
      io_macOut = _22_16_inner_macOut;
    end
  end

  assign _zz__22_16_inner_macOut = ($signed(_zz__zz__22_16_inner_macOut) + $signed(_zz__zz__22_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_16_inner_activation <= 8'h00;
      _22_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_16_inner_activation <= io_addInput;
      end else begin
        _22_16_inner_macOut <= _zz__22_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_719 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_15_inner_macOut;
  wire       [15:0]   _zz__zz__22_15_inner_macOut_1;
  wire       [15:0]   _zz__22_15_inner_macOut_1;
  wire       [15:0]   _zz__22_15_inner_macOut_2;
  reg        [7:0]    _22_15_inner_activation;
  reg        [7:0]    _22_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_15_inner_macOut;

  assign _zz__zz__22_15_inner_macOut = ($signed(io_mulInput) * $signed(_22_15_inner_activation));
  assign _zz__zz__22_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_15_inner_macOut)) ? 16'h007f : _zz__22_15_inner_macOut_2);
  assign _zz__22_15_inner_macOut_2 = (($signed(_zz__22_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_15_inner_activation;
    end else begin
      io_macOut = _22_15_inner_macOut;
    end
  end

  assign _zz__22_15_inner_macOut = ($signed(_zz__zz__22_15_inner_macOut) + $signed(_zz__zz__22_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_15_inner_activation <= 8'h00;
      _22_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_15_inner_activation <= io_addInput;
      end else begin
        _22_15_inner_macOut <= _zz__22_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_718 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_14_inner_macOut;
  wire       [15:0]   _zz__zz__22_14_inner_macOut_1;
  wire       [15:0]   _zz__22_14_inner_macOut_1;
  wire       [15:0]   _zz__22_14_inner_macOut_2;
  reg        [7:0]    _22_14_inner_activation;
  reg        [7:0]    _22_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_14_inner_macOut;

  assign _zz__zz__22_14_inner_macOut = ($signed(io_mulInput) * $signed(_22_14_inner_activation));
  assign _zz__zz__22_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_14_inner_macOut)) ? 16'h007f : _zz__22_14_inner_macOut_2);
  assign _zz__22_14_inner_macOut_2 = (($signed(_zz__22_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_14_inner_activation;
    end else begin
      io_macOut = _22_14_inner_macOut;
    end
  end

  assign _zz__22_14_inner_macOut = ($signed(_zz__zz__22_14_inner_macOut) + $signed(_zz__zz__22_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_14_inner_activation <= 8'h00;
      _22_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_14_inner_activation <= io_addInput;
      end else begin
        _22_14_inner_macOut <= _zz__22_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_717 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_13_inner_macOut;
  wire       [15:0]   _zz__zz__22_13_inner_macOut_1;
  wire       [15:0]   _zz__22_13_inner_macOut_1;
  wire       [15:0]   _zz__22_13_inner_macOut_2;
  reg        [7:0]    _22_13_inner_activation;
  reg        [7:0]    _22_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_13_inner_macOut;

  assign _zz__zz__22_13_inner_macOut = ($signed(io_mulInput) * $signed(_22_13_inner_activation));
  assign _zz__zz__22_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_13_inner_macOut)) ? 16'h007f : _zz__22_13_inner_macOut_2);
  assign _zz__22_13_inner_macOut_2 = (($signed(_zz__22_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_13_inner_activation;
    end else begin
      io_macOut = _22_13_inner_macOut;
    end
  end

  assign _zz__22_13_inner_macOut = ($signed(_zz__zz__22_13_inner_macOut) + $signed(_zz__zz__22_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_13_inner_activation <= 8'h00;
      _22_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_13_inner_activation <= io_addInput;
      end else begin
        _22_13_inner_macOut <= _zz__22_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_716 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_12_inner_macOut;
  wire       [15:0]   _zz__zz__22_12_inner_macOut_1;
  wire       [15:0]   _zz__22_12_inner_macOut_1;
  wire       [15:0]   _zz__22_12_inner_macOut_2;
  reg        [7:0]    _22_12_inner_activation;
  reg        [7:0]    _22_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_12_inner_macOut;

  assign _zz__zz__22_12_inner_macOut = ($signed(io_mulInput) * $signed(_22_12_inner_activation));
  assign _zz__zz__22_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_12_inner_macOut)) ? 16'h007f : _zz__22_12_inner_macOut_2);
  assign _zz__22_12_inner_macOut_2 = (($signed(_zz__22_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_12_inner_activation;
    end else begin
      io_macOut = _22_12_inner_macOut;
    end
  end

  assign _zz__22_12_inner_macOut = ($signed(_zz__zz__22_12_inner_macOut) + $signed(_zz__zz__22_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_12_inner_activation <= 8'h00;
      _22_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_12_inner_activation <= io_addInput;
      end else begin
        _22_12_inner_macOut <= _zz__22_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_715 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_11_inner_macOut;
  wire       [15:0]   _zz__zz__22_11_inner_macOut_1;
  wire       [15:0]   _zz__22_11_inner_macOut_1;
  wire       [15:0]   _zz__22_11_inner_macOut_2;
  reg        [7:0]    _22_11_inner_activation;
  reg        [7:0]    _22_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_11_inner_macOut;

  assign _zz__zz__22_11_inner_macOut = ($signed(io_mulInput) * $signed(_22_11_inner_activation));
  assign _zz__zz__22_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_11_inner_macOut)) ? 16'h007f : _zz__22_11_inner_macOut_2);
  assign _zz__22_11_inner_macOut_2 = (($signed(_zz__22_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_11_inner_activation;
    end else begin
      io_macOut = _22_11_inner_macOut;
    end
  end

  assign _zz__22_11_inner_macOut = ($signed(_zz__zz__22_11_inner_macOut) + $signed(_zz__zz__22_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_11_inner_activation <= 8'h00;
      _22_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_11_inner_activation <= io_addInput;
      end else begin
        _22_11_inner_macOut <= _zz__22_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_714 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_10_inner_macOut;
  wire       [15:0]   _zz__zz__22_10_inner_macOut_1;
  wire       [15:0]   _zz__22_10_inner_macOut_1;
  wire       [15:0]   _zz__22_10_inner_macOut_2;
  reg        [7:0]    _22_10_inner_activation;
  reg        [7:0]    _22_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_10_inner_macOut;

  assign _zz__zz__22_10_inner_macOut = ($signed(io_mulInput) * $signed(_22_10_inner_activation));
  assign _zz__zz__22_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_10_inner_macOut)) ? 16'h007f : _zz__22_10_inner_macOut_2);
  assign _zz__22_10_inner_macOut_2 = (($signed(_zz__22_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_10_inner_activation;
    end else begin
      io_macOut = _22_10_inner_macOut;
    end
  end

  assign _zz__22_10_inner_macOut = ($signed(_zz__zz__22_10_inner_macOut) + $signed(_zz__zz__22_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_10_inner_activation <= 8'h00;
      _22_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_10_inner_activation <= io_addInput;
      end else begin
        _22_10_inner_macOut <= _zz__22_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_713 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_9_inner_macOut;
  wire       [15:0]   _zz__zz__22_9_inner_macOut_1;
  wire       [15:0]   _zz__22_9_inner_macOut_1;
  wire       [15:0]   _zz__22_9_inner_macOut_2;
  reg        [7:0]    _22_9_inner_activation;
  reg        [7:0]    _22_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_9_inner_macOut;

  assign _zz__zz__22_9_inner_macOut = ($signed(io_mulInput) * $signed(_22_9_inner_activation));
  assign _zz__zz__22_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_9_inner_macOut)) ? 16'h007f : _zz__22_9_inner_macOut_2);
  assign _zz__22_9_inner_macOut_2 = (($signed(_zz__22_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_9_inner_activation;
    end else begin
      io_macOut = _22_9_inner_macOut;
    end
  end

  assign _zz__22_9_inner_macOut = ($signed(_zz__zz__22_9_inner_macOut) + $signed(_zz__zz__22_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_9_inner_activation <= 8'h00;
      _22_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_9_inner_activation <= io_addInput;
      end else begin
        _22_9_inner_macOut <= _zz__22_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_712 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_8_inner_macOut;
  wire       [15:0]   _zz__zz__22_8_inner_macOut_1;
  wire       [15:0]   _zz__22_8_inner_macOut_1;
  wire       [15:0]   _zz__22_8_inner_macOut_2;
  reg        [7:0]    _22_8_inner_activation;
  reg        [7:0]    _22_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_8_inner_macOut;

  assign _zz__zz__22_8_inner_macOut = ($signed(io_mulInput) * $signed(_22_8_inner_activation));
  assign _zz__zz__22_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_8_inner_macOut)) ? 16'h007f : _zz__22_8_inner_macOut_2);
  assign _zz__22_8_inner_macOut_2 = (($signed(_zz__22_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_8_inner_activation;
    end else begin
      io_macOut = _22_8_inner_macOut;
    end
  end

  assign _zz__22_8_inner_macOut = ($signed(_zz__zz__22_8_inner_macOut) + $signed(_zz__zz__22_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_8_inner_activation <= 8'h00;
      _22_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_8_inner_activation <= io_addInput;
      end else begin
        _22_8_inner_macOut <= _zz__22_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_711 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_7_inner_macOut;
  wire       [15:0]   _zz__zz__22_7_inner_macOut_1;
  wire       [15:0]   _zz__22_7_inner_macOut_1;
  wire       [15:0]   _zz__22_7_inner_macOut_2;
  reg        [7:0]    _22_7_inner_activation;
  reg        [7:0]    _22_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_7_inner_macOut;

  assign _zz__zz__22_7_inner_macOut = ($signed(io_mulInput) * $signed(_22_7_inner_activation));
  assign _zz__zz__22_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_7_inner_macOut)) ? 16'h007f : _zz__22_7_inner_macOut_2);
  assign _zz__22_7_inner_macOut_2 = (($signed(_zz__22_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_7_inner_activation;
    end else begin
      io_macOut = _22_7_inner_macOut;
    end
  end

  assign _zz__22_7_inner_macOut = ($signed(_zz__zz__22_7_inner_macOut) + $signed(_zz__zz__22_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_7_inner_activation <= 8'h00;
      _22_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_7_inner_activation <= io_addInput;
      end else begin
        _22_7_inner_macOut <= _zz__22_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_710 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_6_inner_macOut;
  wire       [15:0]   _zz__zz__22_6_inner_macOut_1;
  wire       [15:0]   _zz__22_6_inner_macOut_1;
  wire       [15:0]   _zz__22_6_inner_macOut_2;
  reg        [7:0]    _22_6_inner_activation;
  reg        [7:0]    _22_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_6_inner_macOut;

  assign _zz__zz__22_6_inner_macOut = ($signed(io_mulInput) * $signed(_22_6_inner_activation));
  assign _zz__zz__22_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_6_inner_macOut)) ? 16'h007f : _zz__22_6_inner_macOut_2);
  assign _zz__22_6_inner_macOut_2 = (($signed(_zz__22_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_6_inner_activation;
    end else begin
      io_macOut = _22_6_inner_macOut;
    end
  end

  assign _zz__22_6_inner_macOut = ($signed(_zz__zz__22_6_inner_macOut) + $signed(_zz__zz__22_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_6_inner_activation <= 8'h00;
      _22_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_6_inner_activation <= io_addInput;
      end else begin
        _22_6_inner_macOut <= _zz__22_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_709 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_5_inner_macOut;
  wire       [15:0]   _zz__zz__22_5_inner_macOut_1;
  wire       [15:0]   _zz__22_5_inner_macOut_1;
  wire       [15:0]   _zz__22_5_inner_macOut_2;
  reg        [7:0]    _22_5_inner_activation;
  reg        [7:0]    _22_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_5_inner_macOut;

  assign _zz__zz__22_5_inner_macOut = ($signed(io_mulInput) * $signed(_22_5_inner_activation));
  assign _zz__zz__22_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_5_inner_macOut)) ? 16'h007f : _zz__22_5_inner_macOut_2);
  assign _zz__22_5_inner_macOut_2 = (($signed(_zz__22_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_5_inner_activation;
    end else begin
      io_macOut = _22_5_inner_macOut;
    end
  end

  assign _zz__22_5_inner_macOut = ($signed(_zz__zz__22_5_inner_macOut) + $signed(_zz__zz__22_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_5_inner_activation <= 8'h00;
      _22_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_5_inner_activation <= io_addInput;
      end else begin
        _22_5_inner_macOut <= _zz__22_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_708 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_4_inner_macOut;
  wire       [15:0]   _zz__zz__22_4_inner_macOut_1;
  wire       [15:0]   _zz__22_4_inner_macOut_1;
  wire       [15:0]   _zz__22_4_inner_macOut_2;
  reg        [7:0]    _22_4_inner_activation;
  reg        [7:0]    _22_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_4_inner_macOut;

  assign _zz__zz__22_4_inner_macOut = ($signed(io_mulInput) * $signed(_22_4_inner_activation));
  assign _zz__zz__22_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_4_inner_macOut)) ? 16'h007f : _zz__22_4_inner_macOut_2);
  assign _zz__22_4_inner_macOut_2 = (($signed(_zz__22_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_4_inner_activation;
    end else begin
      io_macOut = _22_4_inner_macOut;
    end
  end

  assign _zz__22_4_inner_macOut = ($signed(_zz__zz__22_4_inner_macOut) + $signed(_zz__zz__22_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_4_inner_activation <= 8'h00;
      _22_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_4_inner_activation <= io_addInput;
      end else begin
        _22_4_inner_macOut <= _zz__22_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_707 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_3_inner_macOut;
  wire       [15:0]   _zz__zz__22_3_inner_macOut_1;
  wire       [15:0]   _zz__22_3_inner_macOut_1;
  wire       [15:0]   _zz__22_3_inner_macOut_2;
  reg        [7:0]    _22_3_inner_activation;
  reg        [7:0]    _22_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_3_inner_macOut;

  assign _zz__zz__22_3_inner_macOut = ($signed(io_mulInput) * $signed(_22_3_inner_activation));
  assign _zz__zz__22_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_3_inner_macOut)) ? 16'h007f : _zz__22_3_inner_macOut_2);
  assign _zz__22_3_inner_macOut_2 = (($signed(_zz__22_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_3_inner_activation;
    end else begin
      io_macOut = _22_3_inner_macOut;
    end
  end

  assign _zz__22_3_inner_macOut = ($signed(_zz__zz__22_3_inner_macOut) + $signed(_zz__zz__22_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_3_inner_activation <= 8'h00;
      _22_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_3_inner_activation <= io_addInput;
      end else begin
        _22_3_inner_macOut <= _zz__22_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_706 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_2_inner_macOut;
  wire       [15:0]   _zz__zz__22_2_inner_macOut_1;
  wire       [15:0]   _zz__22_2_inner_macOut_1;
  wire       [15:0]   _zz__22_2_inner_macOut_2;
  reg        [7:0]    _22_2_inner_activation;
  reg        [7:0]    _22_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_2_inner_macOut;

  assign _zz__zz__22_2_inner_macOut = ($signed(io_mulInput) * $signed(_22_2_inner_activation));
  assign _zz__zz__22_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_2_inner_macOut)) ? 16'h007f : _zz__22_2_inner_macOut_2);
  assign _zz__22_2_inner_macOut_2 = (($signed(_zz__22_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_2_inner_activation;
    end else begin
      io_macOut = _22_2_inner_macOut;
    end
  end

  assign _zz__22_2_inner_macOut = ($signed(_zz__zz__22_2_inner_macOut) + $signed(_zz__zz__22_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_2_inner_activation <= 8'h00;
      _22_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_2_inner_activation <= io_addInput;
      end else begin
        _22_2_inner_macOut <= _zz__22_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_705 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_1_inner_macOut;
  wire       [15:0]   _zz__zz__22_1_inner_macOut_1;
  wire       [15:0]   _zz__22_1_inner_macOut_1;
  wire       [15:0]   _zz__22_1_inner_macOut_2;
  reg        [7:0]    _22_1_inner_activation;
  reg        [7:0]    _22_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_1_inner_macOut;

  assign _zz__zz__22_1_inner_macOut = ($signed(io_mulInput) * $signed(_22_1_inner_activation));
  assign _zz__zz__22_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_1_inner_macOut)) ? 16'h007f : _zz__22_1_inner_macOut_2);
  assign _zz__22_1_inner_macOut_2 = (($signed(_zz__22_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_1_inner_activation;
    end else begin
      io_macOut = _22_1_inner_macOut;
    end
  end

  assign _zz__22_1_inner_macOut = ($signed(_zz__zz__22_1_inner_macOut) + $signed(_zz__zz__22_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_1_inner_activation <= 8'h00;
      _22_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_1_inner_activation <= io_addInput;
      end else begin
        _22_1_inner_macOut <= _zz__22_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_704 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__22_0_inner_macOut;
  wire       [15:0]   _zz__zz__22_0_inner_macOut_1;
  wire       [15:0]   _zz__22_0_inner_macOut_1;
  wire       [15:0]   _zz__22_0_inner_macOut_2;
  reg        [7:0]    _22_0_inner_activation;
  reg        [7:0]    _22_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__22_0_inner_macOut;

  assign _zz__zz__22_0_inner_macOut = ($signed(io_mulInput) * $signed(_22_0_inner_activation));
  assign _zz__zz__22_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__22_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__22_0_inner_macOut)) ? 16'h007f : _zz__22_0_inner_macOut_2);
  assign _zz__22_0_inner_macOut_2 = (($signed(_zz__22_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__22_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _22_0_inner_activation;
    end else begin
      io_macOut = _22_0_inner_macOut;
    end
  end

  assign _zz__22_0_inner_macOut = ($signed(_zz__zz__22_0_inner_macOut) + $signed(_zz__zz__22_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _22_0_inner_activation <= 8'h00;
      _22_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _22_0_inner_activation <= io_addInput;
      end else begin
        _22_0_inner_macOut <= _zz__22_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_703 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_31_inner_macOut;
  wire       [15:0]   _zz__zz__21_31_inner_macOut_1;
  wire       [15:0]   _zz__21_31_inner_macOut_1;
  wire       [15:0]   _zz__21_31_inner_macOut_2;
  reg        [7:0]    _21_31_inner_activation;
  reg        [7:0]    _21_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_31_inner_macOut;

  assign _zz__zz__21_31_inner_macOut = ($signed(io_mulInput) * $signed(_21_31_inner_activation));
  assign _zz__zz__21_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_31_inner_macOut)) ? 16'h007f : _zz__21_31_inner_macOut_2);
  assign _zz__21_31_inner_macOut_2 = (($signed(_zz__21_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_31_inner_activation;
    end else begin
      io_macOut = _21_31_inner_macOut;
    end
  end

  assign _zz__21_31_inner_macOut = ($signed(_zz__zz__21_31_inner_macOut) + $signed(_zz__zz__21_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_31_inner_activation <= 8'h00;
      _21_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_31_inner_activation <= io_addInput;
      end else begin
        _21_31_inner_macOut <= _zz__21_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_702 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_30_inner_macOut;
  wire       [15:0]   _zz__zz__21_30_inner_macOut_1;
  wire       [15:0]   _zz__21_30_inner_macOut_1;
  wire       [15:0]   _zz__21_30_inner_macOut_2;
  reg        [7:0]    _21_30_inner_activation;
  reg        [7:0]    _21_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_30_inner_macOut;

  assign _zz__zz__21_30_inner_macOut = ($signed(io_mulInput) * $signed(_21_30_inner_activation));
  assign _zz__zz__21_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_30_inner_macOut)) ? 16'h007f : _zz__21_30_inner_macOut_2);
  assign _zz__21_30_inner_macOut_2 = (($signed(_zz__21_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_30_inner_activation;
    end else begin
      io_macOut = _21_30_inner_macOut;
    end
  end

  assign _zz__21_30_inner_macOut = ($signed(_zz__zz__21_30_inner_macOut) + $signed(_zz__zz__21_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_30_inner_activation <= 8'h00;
      _21_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_30_inner_activation <= io_addInput;
      end else begin
        _21_30_inner_macOut <= _zz__21_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_701 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_29_inner_macOut;
  wire       [15:0]   _zz__zz__21_29_inner_macOut_1;
  wire       [15:0]   _zz__21_29_inner_macOut_1;
  wire       [15:0]   _zz__21_29_inner_macOut_2;
  reg        [7:0]    _21_29_inner_activation;
  reg        [7:0]    _21_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_29_inner_macOut;

  assign _zz__zz__21_29_inner_macOut = ($signed(io_mulInput) * $signed(_21_29_inner_activation));
  assign _zz__zz__21_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_29_inner_macOut)) ? 16'h007f : _zz__21_29_inner_macOut_2);
  assign _zz__21_29_inner_macOut_2 = (($signed(_zz__21_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_29_inner_activation;
    end else begin
      io_macOut = _21_29_inner_macOut;
    end
  end

  assign _zz__21_29_inner_macOut = ($signed(_zz__zz__21_29_inner_macOut) + $signed(_zz__zz__21_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_29_inner_activation <= 8'h00;
      _21_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_29_inner_activation <= io_addInput;
      end else begin
        _21_29_inner_macOut <= _zz__21_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_700 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_28_inner_macOut;
  wire       [15:0]   _zz__zz__21_28_inner_macOut_1;
  wire       [15:0]   _zz__21_28_inner_macOut_1;
  wire       [15:0]   _zz__21_28_inner_macOut_2;
  reg        [7:0]    _21_28_inner_activation;
  reg        [7:0]    _21_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_28_inner_macOut;

  assign _zz__zz__21_28_inner_macOut = ($signed(io_mulInput) * $signed(_21_28_inner_activation));
  assign _zz__zz__21_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_28_inner_macOut)) ? 16'h007f : _zz__21_28_inner_macOut_2);
  assign _zz__21_28_inner_macOut_2 = (($signed(_zz__21_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_28_inner_activation;
    end else begin
      io_macOut = _21_28_inner_macOut;
    end
  end

  assign _zz__21_28_inner_macOut = ($signed(_zz__zz__21_28_inner_macOut) + $signed(_zz__zz__21_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_28_inner_activation <= 8'h00;
      _21_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_28_inner_activation <= io_addInput;
      end else begin
        _21_28_inner_macOut <= _zz__21_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_699 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_27_inner_macOut;
  wire       [15:0]   _zz__zz__21_27_inner_macOut_1;
  wire       [15:0]   _zz__21_27_inner_macOut_1;
  wire       [15:0]   _zz__21_27_inner_macOut_2;
  reg        [7:0]    _21_27_inner_activation;
  reg        [7:0]    _21_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_27_inner_macOut;

  assign _zz__zz__21_27_inner_macOut = ($signed(io_mulInput) * $signed(_21_27_inner_activation));
  assign _zz__zz__21_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_27_inner_macOut)) ? 16'h007f : _zz__21_27_inner_macOut_2);
  assign _zz__21_27_inner_macOut_2 = (($signed(_zz__21_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_27_inner_activation;
    end else begin
      io_macOut = _21_27_inner_macOut;
    end
  end

  assign _zz__21_27_inner_macOut = ($signed(_zz__zz__21_27_inner_macOut) + $signed(_zz__zz__21_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_27_inner_activation <= 8'h00;
      _21_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_27_inner_activation <= io_addInput;
      end else begin
        _21_27_inner_macOut <= _zz__21_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_698 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_26_inner_macOut;
  wire       [15:0]   _zz__zz__21_26_inner_macOut_1;
  wire       [15:0]   _zz__21_26_inner_macOut_1;
  wire       [15:0]   _zz__21_26_inner_macOut_2;
  reg        [7:0]    _21_26_inner_activation;
  reg        [7:0]    _21_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_26_inner_macOut;

  assign _zz__zz__21_26_inner_macOut = ($signed(io_mulInput) * $signed(_21_26_inner_activation));
  assign _zz__zz__21_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_26_inner_macOut)) ? 16'h007f : _zz__21_26_inner_macOut_2);
  assign _zz__21_26_inner_macOut_2 = (($signed(_zz__21_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_26_inner_activation;
    end else begin
      io_macOut = _21_26_inner_macOut;
    end
  end

  assign _zz__21_26_inner_macOut = ($signed(_zz__zz__21_26_inner_macOut) + $signed(_zz__zz__21_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_26_inner_activation <= 8'h00;
      _21_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_26_inner_activation <= io_addInput;
      end else begin
        _21_26_inner_macOut <= _zz__21_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_697 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_25_inner_macOut;
  wire       [15:0]   _zz__zz__21_25_inner_macOut_1;
  wire       [15:0]   _zz__21_25_inner_macOut_1;
  wire       [15:0]   _zz__21_25_inner_macOut_2;
  reg        [7:0]    _21_25_inner_activation;
  reg        [7:0]    _21_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_25_inner_macOut;

  assign _zz__zz__21_25_inner_macOut = ($signed(io_mulInput) * $signed(_21_25_inner_activation));
  assign _zz__zz__21_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_25_inner_macOut)) ? 16'h007f : _zz__21_25_inner_macOut_2);
  assign _zz__21_25_inner_macOut_2 = (($signed(_zz__21_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_25_inner_activation;
    end else begin
      io_macOut = _21_25_inner_macOut;
    end
  end

  assign _zz__21_25_inner_macOut = ($signed(_zz__zz__21_25_inner_macOut) + $signed(_zz__zz__21_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_25_inner_activation <= 8'h00;
      _21_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_25_inner_activation <= io_addInput;
      end else begin
        _21_25_inner_macOut <= _zz__21_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_696 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_24_inner_macOut;
  wire       [15:0]   _zz__zz__21_24_inner_macOut_1;
  wire       [15:0]   _zz__21_24_inner_macOut_1;
  wire       [15:0]   _zz__21_24_inner_macOut_2;
  reg        [7:0]    _21_24_inner_activation;
  reg        [7:0]    _21_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_24_inner_macOut;

  assign _zz__zz__21_24_inner_macOut = ($signed(io_mulInput) * $signed(_21_24_inner_activation));
  assign _zz__zz__21_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_24_inner_macOut)) ? 16'h007f : _zz__21_24_inner_macOut_2);
  assign _zz__21_24_inner_macOut_2 = (($signed(_zz__21_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_24_inner_activation;
    end else begin
      io_macOut = _21_24_inner_macOut;
    end
  end

  assign _zz__21_24_inner_macOut = ($signed(_zz__zz__21_24_inner_macOut) + $signed(_zz__zz__21_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_24_inner_activation <= 8'h00;
      _21_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_24_inner_activation <= io_addInput;
      end else begin
        _21_24_inner_macOut <= _zz__21_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_695 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_23_inner_macOut;
  wire       [15:0]   _zz__zz__21_23_inner_macOut_1;
  wire       [15:0]   _zz__21_23_inner_macOut_1;
  wire       [15:0]   _zz__21_23_inner_macOut_2;
  reg        [7:0]    _21_23_inner_activation;
  reg        [7:0]    _21_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_23_inner_macOut;

  assign _zz__zz__21_23_inner_macOut = ($signed(io_mulInput) * $signed(_21_23_inner_activation));
  assign _zz__zz__21_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_23_inner_macOut)) ? 16'h007f : _zz__21_23_inner_macOut_2);
  assign _zz__21_23_inner_macOut_2 = (($signed(_zz__21_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_23_inner_activation;
    end else begin
      io_macOut = _21_23_inner_macOut;
    end
  end

  assign _zz__21_23_inner_macOut = ($signed(_zz__zz__21_23_inner_macOut) + $signed(_zz__zz__21_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_23_inner_activation <= 8'h00;
      _21_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_23_inner_activation <= io_addInput;
      end else begin
        _21_23_inner_macOut <= _zz__21_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_694 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_22_inner_macOut;
  wire       [15:0]   _zz__zz__21_22_inner_macOut_1;
  wire       [15:0]   _zz__21_22_inner_macOut_1;
  wire       [15:0]   _zz__21_22_inner_macOut_2;
  reg        [7:0]    _21_22_inner_activation;
  reg        [7:0]    _21_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_22_inner_macOut;

  assign _zz__zz__21_22_inner_macOut = ($signed(io_mulInput) * $signed(_21_22_inner_activation));
  assign _zz__zz__21_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_22_inner_macOut)) ? 16'h007f : _zz__21_22_inner_macOut_2);
  assign _zz__21_22_inner_macOut_2 = (($signed(_zz__21_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_22_inner_activation;
    end else begin
      io_macOut = _21_22_inner_macOut;
    end
  end

  assign _zz__21_22_inner_macOut = ($signed(_zz__zz__21_22_inner_macOut) + $signed(_zz__zz__21_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_22_inner_activation <= 8'h00;
      _21_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_22_inner_activation <= io_addInput;
      end else begin
        _21_22_inner_macOut <= _zz__21_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_693 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_21_inner_macOut;
  wire       [15:0]   _zz__zz__21_21_inner_macOut_1;
  wire       [15:0]   _zz__21_21_inner_macOut_1;
  wire       [15:0]   _zz__21_21_inner_macOut_2;
  reg        [7:0]    _21_21_inner_activation;
  reg        [7:0]    _21_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_21_inner_macOut;

  assign _zz__zz__21_21_inner_macOut = ($signed(io_mulInput) * $signed(_21_21_inner_activation));
  assign _zz__zz__21_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_21_inner_macOut)) ? 16'h007f : _zz__21_21_inner_macOut_2);
  assign _zz__21_21_inner_macOut_2 = (($signed(_zz__21_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_21_inner_activation;
    end else begin
      io_macOut = _21_21_inner_macOut;
    end
  end

  assign _zz__21_21_inner_macOut = ($signed(_zz__zz__21_21_inner_macOut) + $signed(_zz__zz__21_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_21_inner_activation <= 8'h00;
      _21_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_21_inner_activation <= io_addInput;
      end else begin
        _21_21_inner_macOut <= _zz__21_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_692 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_20_inner_macOut;
  wire       [15:0]   _zz__zz__21_20_inner_macOut_1;
  wire       [15:0]   _zz__21_20_inner_macOut_1;
  wire       [15:0]   _zz__21_20_inner_macOut_2;
  reg        [7:0]    _21_20_inner_activation;
  reg        [7:0]    _21_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_20_inner_macOut;

  assign _zz__zz__21_20_inner_macOut = ($signed(io_mulInput) * $signed(_21_20_inner_activation));
  assign _zz__zz__21_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_20_inner_macOut)) ? 16'h007f : _zz__21_20_inner_macOut_2);
  assign _zz__21_20_inner_macOut_2 = (($signed(_zz__21_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_20_inner_activation;
    end else begin
      io_macOut = _21_20_inner_macOut;
    end
  end

  assign _zz__21_20_inner_macOut = ($signed(_zz__zz__21_20_inner_macOut) + $signed(_zz__zz__21_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_20_inner_activation <= 8'h00;
      _21_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_20_inner_activation <= io_addInput;
      end else begin
        _21_20_inner_macOut <= _zz__21_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_691 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_19_inner_macOut;
  wire       [15:0]   _zz__zz__21_19_inner_macOut_1;
  wire       [15:0]   _zz__21_19_inner_macOut_1;
  wire       [15:0]   _zz__21_19_inner_macOut_2;
  reg        [7:0]    _21_19_inner_activation;
  reg        [7:0]    _21_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_19_inner_macOut;

  assign _zz__zz__21_19_inner_macOut = ($signed(io_mulInput) * $signed(_21_19_inner_activation));
  assign _zz__zz__21_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_19_inner_macOut)) ? 16'h007f : _zz__21_19_inner_macOut_2);
  assign _zz__21_19_inner_macOut_2 = (($signed(_zz__21_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_19_inner_activation;
    end else begin
      io_macOut = _21_19_inner_macOut;
    end
  end

  assign _zz__21_19_inner_macOut = ($signed(_zz__zz__21_19_inner_macOut) + $signed(_zz__zz__21_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_19_inner_activation <= 8'h00;
      _21_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_19_inner_activation <= io_addInput;
      end else begin
        _21_19_inner_macOut <= _zz__21_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_690 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_18_inner_macOut;
  wire       [15:0]   _zz__zz__21_18_inner_macOut_1;
  wire       [15:0]   _zz__21_18_inner_macOut_1;
  wire       [15:0]   _zz__21_18_inner_macOut_2;
  reg        [7:0]    _21_18_inner_activation;
  reg        [7:0]    _21_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_18_inner_macOut;

  assign _zz__zz__21_18_inner_macOut = ($signed(io_mulInput) * $signed(_21_18_inner_activation));
  assign _zz__zz__21_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_18_inner_macOut)) ? 16'h007f : _zz__21_18_inner_macOut_2);
  assign _zz__21_18_inner_macOut_2 = (($signed(_zz__21_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_18_inner_activation;
    end else begin
      io_macOut = _21_18_inner_macOut;
    end
  end

  assign _zz__21_18_inner_macOut = ($signed(_zz__zz__21_18_inner_macOut) + $signed(_zz__zz__21_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_18_inner_activation <= 8'h00;
      _21_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_18_inner_activation <= io_addInput;
      end else begin
        _21_18_inner_macOut <= _zz__21_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_689 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_17_inner_macOut;
  wire       [15:0]   _zz__zz__21_17_inner_macOut_1;
  wire       [15:0]   _zz__21_17_inner_macOut_1;
  wire       [15:0]   _zz__21_17_inner_macOut_2;
  reg        [7:0]    _21_17_inner_activation;
  reg        [7:0]    _21_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_17_inner_macOut;

  assign _zz__zz__21_17_inner_macOut = ($signed(io_mulInput) * $signed(_21_17_inner_activation));
  assign _zz__zz__21_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_17_inner_macOut)) ? 16'h007f : _zz__21_17_inner_macOut_2);
  assign _zz__21_17_inner_macOut_2 = (($signed(_zz__21_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_17_inner_activation;
    end else begin
      io_macOut = _21_17_inner_macOut;
    end
  end

  assign _zz__21_17_inner_macOut = ($signed(_zz__zz__21_17_inner_macOut) + $signed(_zz__zz__21_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_17_inner_activation <= 8'h00;
      _21_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_17_inner_activation <= io_addInput;
      end else begin
        _21_17_inner_macOut <= _zz__21_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_688 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_16_inner_macOut;
  wire       [15:0]   _zz__zz__21_16_inner_macOut_1;
  wire       [15:0]   _zz__21_16_inner_macOut_1;
  wire       [15:0]   _zz__21_16_inner_macOut_2;
  reg        [7:0]    _21_16_inner_activation;
  reg        [7:0]    _21_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_16_inner_macOut;

  assign _zz__zz__21_16_inner_macOut = ($signed(io_mulInput) * $signed(_21_16_inner_activation));
  assign _zz__zz__21_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_16_inner_macOut)) ? 16'h007f : _zz__21_16_inner_macOut_2);
  assign _zz__21_16_inner_macOut_2 = (($signed(_zz__21_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_16_inner_activation;
    end else begin
      io_macOut = _21_16_inner_macOut;
    end
  end

  assign _zz__21_16_inner_macOut = ($signed(_zz__zz__21_16_inner_macOut) + $signed(_zz__zz__21_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_16_inner_activation <= 8'h00;
      _21_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_16_inner_activation <= io_addInput;
      end else begin
        _21_16_inner_macOut <= _zz__21_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_687 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_15_inner_macOut;
  wire       [15:0]   _zz__zz__21_15_inner_macOut_1;
  wire       [15:0]   _zz__21_15_inner_macOut_1;
  wire       [15:0]   _zz__21_15_inner_macOut_2;
  reg        [7:0]    _21_15_inner_activation;
  reg        [7:0]    _21_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_15_inner_macOut;

  assign _zz__zz__21_15_inner_macOut = ($signed(io_mulInput) * $signed(_21_15_inner_activation));
  assign _zz__zz__21_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_15_inner_macOut)) ? 16'h007f : _zz__21_15_inner_macOut_2);
  assign _zz__21_15_inner_macOut_2 = (($signed(_zz__21_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_15_inner_activation;
    end else begin
      io_macOut = _21_15_inner_macOut;
    end
  end

  assign _zz__21_15_inner_macOut = ($signed(_zz__zz__21_15_inner_macOut) + $signed(_zz__zz__21_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_15_inner_activation <= 8'h00;
      _21_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_15_inner_activation <= io_addInput;
      end else begin
        _21_15_inner_macOut <= _zz__21_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_686 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_14_inner_macOut;
  wire       [15:0]   _zz__zz__21_14_inner_macOut_1;
  wire       [15:0]   _zz__21_14_inner_macOut_1;
  wire       [15:0]   _zz__21_14_inner_macOut_2;
  reg        [7:0]    _21_14_inner_activation;
  reg        [7:0]    _21_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_14_inner_macOut;

  assign _zz__zz__21_14_inner_macOut = ($signed(io_mulInput) * $signed(_21_14_inner_activation));
  assign _zz__zz__21_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_14_inner_macOut)) ? 16'h007f : _zz__21_14_inner_macOut_2);
  assign _zz__21_14_inner_macOut_2 = (($signed(_zz__21_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_14_inner_activation;
    end else begin
      io_macOut = _21_14_inner_macOut;
    end
  end

  assign _zz__21_14_inner_macOut = ($signed(_zz__zz__21_14_inner_macOut) + $signed(_zz__zz__21_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_14_inner_activation <= 8'h00;
      _21_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_14_inner_activation <= io_addInput;
      end else begin
        _21_14_inner_macOut <= _zz__21_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_685 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_13_inner_macOut;
  wire       [15:0]   _zz__zz__21_13_inner_macOut_1;
  wire       [15:0]   _zz__21_13_inner_macOut_1;
  wire       [15:0]   _zz__21_13_inner_macOut_2;
  reg        [7:0]    _21_13_inner_activation;
  reg        [7:0]    _21_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_13_inner_macOut;

  assign _zz__zz__21_13_inner_macOut = ($signed(io_mulInput) * $signed(_21_13_inner_activation));
  assign _zz__zz__21_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_13_inner_macOut)) ? 16'h007f : _zz__21_13_inner_macOut_2);
  assign _zz__21_13_inner_macOut_2 = (($signed(_zz__21_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_13_inner_activation;
    end else begin
      io_macOut = _21_13_inner_macOut;
    end
  end

  assign _zz__21_13_inner_macOut = ($signed(_zz__zz__21_13_inner_macOut) + $signed(_zz__zz__21_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_13_inner_activation <= 8'h00;
      _21_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_13_inner_activation <= io_addInput;
      end else begin
        _21_13_inner_macOut <= _zz__21_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_684 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_12_inner_macOut;
  wire       [15:0]   _zz__zz__21_12_inner_macOut_1;
  wire       [15:0]   _zz__21_12_inner_macOut_1;
  wire       [15:0]   _zz__21_12_inner_macOut_2;
  reg        [7:0]    _21_12_inner_activation;
  reg        [7:0]    _21_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_12_inner_macOut;

  assign _zz__zz__21_12_inner_macOut = ($signed(io_mulInput) * $signed(_21_12_inner_activation));
  assign _zz__zz__21_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_12_inner_macOut)) ? 16'h007f : _zz__21_12_inner_macOut_2);
  assign _zz__21_12_inner_macOut_2 = (($signed(_zz__21_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_12_inner_activation;
    end else begin
      io_macOut = _21_12_inner_macOut;
    end
  end

  assign _zz__21_12_inner_macOut = ($signed(_zz__zz__21_12_inner_macOut) + $signed(_zz__zz__21_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_12_inner_activation <= 8'h00;
      _21_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_12_inner_activation <= io_addInput;
      end else begin
        _21_12_inner_macOut <= _zz__21_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_683 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_11_inner_macOut;
  wire       [15:0]   _zz__zz__21_11_inner_macOut_1;
  wire       [15:0]   _zz__21_11_inner_macOut_1;
  wire       [15:0]   _zz__21_11_inner_macOut_2;
  reg        [7:0]    _21_11_inner_activation;
  reg        [7:0]    _21_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_11_inner_macOut;

  assign _zz__zz__21_11_inner_macOut = ($signed(io_mulInput) * $signed(_21_11_inner_activation));
  assign _zz__zz__21_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_11_inner_macOut)) ? 16'h007f : _zz__21_11_inner_macOut_2);
  assign _zz__21_11_inner_macOut_2 = (($signed(_zz__21_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_11_inner_activation;
    end else begin
      io_macOut = _21_11_inner_macOut;
    end
  end

  assign _zz__21_11_inner_macOut = ($signed(_zz__zz__21_11_inner_macOut) + $signed(_zz__zz__21_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_11_inner_activation <= 8'h00;
      _21_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_11_inner_activation <= io_addInput;
      end else begin
        _21_11_inner_macOut <= _zz__21_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_682 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_10_inner_macOut;
  wire       [15:0]   _zz__zz__21_10_inner_macOut_1;
  wire       [15:0]   _zz__21_10_inner_macOut_1;
  wire       [15:0]   _zz__21_10_inner_macOut_2;
  reg        [7:0]    _21_10_inner_activation;
  reg        [7:0]    _21_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_10_inner_macOut;

  assign _zz__zz__21_10_inner_macOut = ($signed(io_mulInput) * $signed(_21_10_inner_activation));
  assign _zz__zz__21_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_10_inner_macOut)) ? 16'h007f : _zz__21_10_inner_macOut_2);
  assign _zz__21_10_inner_macOut_2 = (($signed(_zz__21_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_10_inner_activation;
    end else begin
      io_macOut = _21_10_inner_macOut;
    end
  end

  assign _zz__21_10_inner_macOut = ($signed(_zz__zz__21_10_inner_macOut) + $signed(_zz__zz__21_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_10_inner_activation <= 8'h00;
      _21_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_10_inner_activation <= io_addInput;
      end else begin
        _21_10_inner_macOut <= _zz__21_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_681 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_9_inner_macOut;
  wire       [15:0]   _zz__zz__21_9_inner_macOut_1;
  wire       [15:0]   _zz__21_9_inner_macOut_1;
  wire       [15:0]   _zz__21_9_inner_macOut_2;
  reg        [7:0]    _21_9_inner_activation;
  reg        [7:0]    _21_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_9_inner_macOut;

  assign _zz__zz__21_9_inner_macOut = ($signed(io_mulInput) * $signed(_21_9_inner_activation));
  assign _zz__zz__21_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_9_inner_macOut)) ? 16'h007f : _zz__21_9_inner_macOut_2);
  assign _zz__21_9_inner_macOut_2 = (($signed(_zz__21_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_9_inner_activation;
    end else begin
      io_macOut = _21_9_inner_macOut;
    end
  end

  assign _zz__21_9_inner_macOut = ($signed(_zz__zz__21_9_inner_macOut) + $signed(_zz__zz__21_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_9_inner_activation <= 8'h00;
      _21_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_9_inner_activation <= io_addInput;
      end else begin
        _21_9_inner_macOut <= _zz__21_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_680 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_8_inner_macOut;
  wire       [15:0]   _zz__zz__21_8_inner_macOut_1;
  wire       [15:0]   _zz__21_8_inner_macOut_1;
  wire       [15:0]   _zz__21_8_inner_macOut_2;
  reg        [7:0]    _21_8_inner_activation;
  reg        [7:0]    _21_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_8_inner_macOut;

  assign _zz__zz__21_8_inner_macOut = ($signed(io_mulInput) * $signed(_21_8_inner_activation));
  assign _zz__zz__21_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_8_inner_macOut)) ? 16'h007f : _zz__21_8_inner_macOut_2);
  assign _zz__21_8_inner_macOut_2 = (($signed(_zz__21_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_8_inner_activation;
    end else begin
      io_macOut = _21_8_inner_macOut;
    end
  end

  assign _zz__21_8_inner_macOut = ($signed(_zz__zz__21_8_inner_macOut) + $signed(_zz__zz__21_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_8_inner_activation <= 8'h00;
      _21_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_8_inner_activation <= io_addInput;
      end else begin
        _21_8_inner_macOut <= _zz__21_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_679 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_7_inner_macOut;
  wire       [15:0]   _zz__zz__21_7_inner_macOut_1;
  wire       [15:0]   _zz__21_7_inner_macOut_1;
  wire       [15:0]   _zz__21_7_inner_macOut_2;
  reg        [7:0]    _21_7_inner_activation;
  reg        [7:0]    _21_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_7_inner_macOut;

  assign _zz__zz__21_7_inner_macOut = ($signed(io_mulInput) * $signed(_21_7_inner_activation));
  assign _zz__zz__21_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_7_inner_macOut)) ? 16'h007f : _zz__21_7_inner_macOut_2);
  assign _zz__21_7_inner_macOut_2 = (($signed(_zz__21_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_7_inner_activation;
    end else begin
      io_macOut = _21_7_inner_macOut;
    end
  end

  assign _zz__21_7_inner_macOut = ($signed(_zz__zz__21_7_inner_macOut) + $signed(_zz__zz__21_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_7_inner_activation <= 8'h00;
      _21_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_7_inner_activation <= io_addInput;
      end else begin
        _21_7_inner_macOut <= _zz__21_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_678 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_6_inner_macOut;
  wire       [15:0]   _zz__zz__21_6_inner_macOut_1;
  wire       [15:0]   _zz__21_6_inner_macOut_1;
  wire       [15:0]   _zz__21_6_inner_macOut_2;
  reg        [7:0]    _21_6_inner_activation;
  reg        [7:0]    _21_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_6_inner_macOut;

  assign _zz__zz__21_6_inner_macOut = ($signed(io_mulInput) * $signed(_21_6_inner_activation));
  assign _zz__zz__21_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_6_inner_macOut)) ? 16'h007f : _zz__21_6_inner_macOut_2);
  assign _zz__21_6_inner_macOut_2 = (($signed(_zz__21_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_6_inner_activation;
    end else begin
      io_macOut = _21_6_inner_macOut;
    end
  end

  assign _zz__21_6_inner_macOut = ($signed(_zz__zz__21_6_inner_macOut) + $signed(_zz__zz__21_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_6_inner_activation <= 8'h00;
      _21_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_6_inner_activation <= io_addInput;
      end else begin
        _21_6_inner_macOut <= _zz__21_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_677 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_5_inner_macOut;
  wire       [15:0]   _zz__zz__21_5_inner_macOut_1;
  wire       [15:0]   _zz__21_5_inner_macOut_1;
  wire       [15:0]   _zz__21_5_inner_macOut_2;
  reg        [7:0]    _21_5_inner_activation;
  reg        [7:0]    _21_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_5_inner_macOut;

  assign _zz__zz__21_5_inner_macOut = ($signed(io_mulInput) * $signed(_21_5_inner_activation));
  assign _zz__zz__21_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_5_inner_macOut)) ? 16'h007f : _zz__21_5_inner_macOut_2);
  assign _zz__21_5_inner_macOut_2 = (($signed(_zz__21_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_5_inner_activation;
    end else begin
      io_macOut = _21_5_inner_macOut;
    end
  end

  assign _zz__21_5_inner_macOut = ($signed(_zz__zz__21_5_inner_macOut) + $signed(_zz__zz__21_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_5_inner_activation <= 8'h00;
      _21_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_5_inner_activation <= io_addInput;
      end else begin
        _21_5_inner_macOut <= _zz__21_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_676 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_4_inner_macOut;
  wire       [15:0]   _zz__zz__21_4_inner_macOut_1;
  wire       [15:0]   _zz__21_4_inner_macOut_1;
  wire       [15:0]   _zz__21_4_inner_macOut_2;
  reg        [7:0]    _21_4_inner_activation;
  reg        [7:0]    _21_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_4_inner_macOut;

  assign _zz__zz__21_4_inner_macOut = ($signed(io_mulInput) * $signed(_21_4_inner_activation));
  assign _zz__zz__21_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_4_inner_macOut)) ? 16'h007f : _zz__21_4_inner_macOut_2);
  assign _zz__21_4_inner_macOut_2 = (($signed(_zz__21_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_4_inner_activation;
    end else begin
      io_macOut = _21_4_inner_macOut;
    end
  end

  assign _zz__21_4_inner_macOut = ($signed(_zz__zz__21_4_inner_macOut) + $signed(_zz__zz__21_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_4_inner_activation <= 8'h00;
      _21_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_4_inner_activation <= io_addInput;
      end else begin
        _21_4_inner_macOut <= _zz__21_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_675 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_3_inner_macOut;
  wire       [15:0]   _zz__zz__21_3_inner_macOut_1;
  wire       [15:0]   _zz__21_3_inner_macOut_1;
  wire       [15:0]   _zz__21_3_inner_macOut_2;
  reg        [7:0]    _21_3_inner_activation;
  reg        [7:0]    _21_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_3_inner_macOut;

  assign _zz__zz__21_3_inner_macOut = ($signed(io_mulInput) * $signed(_21_3_inner_activation));
  assign _zz__zz__21_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_3_inner_macOut)) ? 16'h007f : _zz__21_3_inner_macOut_2);
  assign _zz__21_3_inner_macOut_2 = (($signed(_zz__21_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_3_inner_activation;
    end else begin
      io_macOut = _21_3_inner_macOut;
    end
  end

  assign _zz__21_3_inner_macOut = ($signed(_zz__zz__21_3_inner_macOut) + $signed(_zz__zz__21_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_3_inner_activation <= 8'h00;
      _21_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_3_inner_activation <= io_addInput;
      end else begin
        _21_3_inner_macOut <= _zz__21_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_674 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_2_inner_macOut;
  wire       [15:0]   _zz__zz__21_2_inner_macOut_1;
  wire       [15:0]   _zz__21_2_inner_macOut_1;
  wire       [15:0]   _zz__21_2_inner_macOut_2;
  reg        [7:0]    _21_2_inner_activation;
  reg        [7:0]    _21_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_2_inner_macOut;

  assign _zz__zz__21_2_inner_macOut = ($signed(io_mulInput) * $signed(_21_2_inner_activation));
  assign _zz__zz__21_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_2_inner_macOut)) ? 16'h007f : _zz__21_2_inner_macOut_2);
  assign _zz__21_2_inner_macOut_2 = (($signed(_zz__21_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_2_inner_activation;
    end else begin
      io_macOut = _21_2_inner_macOut;
    end
  end

  assign _zz__21_2_inner_macOut = ($signed(_zz__zz__21_2_inner_macOut) + $signed(_zz__zz__21_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_2_inner_activation <= 8'h00;
      _21_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_2_inner_activation <= io_addInput;
      end else begin
        _21_2_inner_macOut <= _zz__21_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_673 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_1_inner_macOut;
  wire       [15:0]   _zz__zz__21_1_inner_macOut_1;
  wire       [15:0]   _zz__21_1_inner_macOut_1;
  wire       [15:0]   _zz__21_1_inner_macOut_2;
  reg        [7:0]    _21_1_inner_activation;
  reg        [7:0]    _21_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_1_inner_macOut;

  assign _zz__zz__21_1_inner_macOut = ($signed(io_mulInput) * $signed(_21_1_inner_activation));
  assign _zz__zz__21_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_1_inner_macOut)) ? 16'h007f : _zz__21_1_inner_macOut_2);
  assign _zz__21_1_inner_macOut_2 = (($signed(_zz__21_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_1_inner_activation;
    end else begin
      io_macOut = _21_1_inner_macOut;
    end
  end

  assign _zz__21_1_inner_macOut = ($signed(_zz__zz__21_1_inner_macOut) + $signed(_zz__zz__21_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_1_inner_activation <= 8'h00;
      _21_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_1_inner_activation <= io_addInput;
      end else begin
        _21_1_inner_macOut <= _zz__21_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_672 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__21_0_inner_macOut;
  wire       [15:0]   _zz__zz__21_0_inner_macOut_1;
  wire       [15:0]   _zz__21_0_inner_macOut_1;
  wire       [15:0]   _zz__21_0_inner_macOut_2;
  reg        [7:0]    _21_0_inner_activation;
  reg        [7:0]    _21_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__21_0_inner_macOut;

  assign _zz__zz__21_0_inner_macOut = ($signed(io_mulInput) * $signed(_21_0_inner_activation));
  assign _zz__zz__21_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__21_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__21_0_inner_macOut)) ? 16'h007f : _zz__21_0_inner_macOut_2);
  assign _zz__21_0_inner_macOut_2 = (($signed(_zz__21_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__21_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _21_0_inner_activation;
    end else begin
      io_macOut = _21_0_inner_macOut;
    end
  end

  assign _zz__21_0_inner_macOut = ($signed(_zz__zz__21_0_inner_macOut) + $signed(_zz__zz__21_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _21_0_inner_activation <= 8'h00;
      _21_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _21_0_inner_activation <= io_addInput;
      end else begin
        _21_0_inner_macOut <= _zz__21_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_671 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_31_inner_macOut;
  wire       [15:0]   _zz__zz__20_31_inner_macOut_1;
  wire       [15:0]   _zz__20_31_inner_macOut_1;
  wire       [15:0]   _zz__20_31_inner_macOut_2;
  reg        [7:0]    _20_31_inner_activation;
  reg        [7:0]    _20_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_31_inner_macOut;

  assign _zz__zz__20_31_inner_macOut = ($signed(io_mulInput) * $signed(_20_31_inner_activation));
  assign _zz__zz__20_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_31_inner_macOut)) ? 16'h007f : _zz__20_31_inner_macOut_2);
  assign _zz__20_31_inner_macOut_2 = (($signed(_zz__20_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_31_inner_activation;
    end else begin
      io_macOut = _20_31_inner_macOut;
    end
  end

  assign _zz__20_31_inner_macOut = ($signed(_zz__zz__20_31_inner_macOut) + $signed(_zz__zz__20_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_31_inner_activation <= 8'h00;
      _20_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_31_inner_activation <= io_addInput;
      end else begin
        _20_31_inner_macOut <= _zz__20_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_670 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_30_inner_macOut;
  wire       [15:0]   _zz__zz__20_30_inner_macOut_1;
  wire       [15:0]   _zz__20_30_inner_macOut_1;
  wire       [15:0]   _zz__20_30_inner_macOut_2;
  reg        [7:0]    _20_30_inner_activation;
  reg        [7:0]    _20_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_30_inner_macOut;

  assign _zz__zz__20_30_inner_macOut = ($signed(io_mulInput) * $signed(_20_30_inner_activation));
  assign _zz__zz__20_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_30_inner_macOut)) ? 16'h007f : _zz__20_30_inner_macOut_2);
  assign _zz__20_30_inner_macOut_2 = (($signed(_zz__20_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_30_inner_activation;
    end else begin
      io_macOut = _20_30_inner_macOut;
    end
  end

  assign _zz__20_30_inner_macOut = ($signed(_zz__zz__20_30_inner_macOut) + $signed(_zz__zz__20_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_30_inner_activation <= 8'h00;
      _20_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_30_inner_activation <= io_addInput;
      end else begin
        _20_30_inner_macOut <= _zz__20_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_669 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_29_inner_macOut;
  wire       [15:0]   _zz__zz__20_29_inner_macOut_1;
  wire       [15:0]   _zz__20_29_inner_macOut_1;
  wire       [15:0]   _zz__20_29_inner_macOut_2;
  reg        [7:0]    _20_29_inner_activation;
  reg        [7:0]    _20_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_29_inner_macOut;

  assign _zz__zz__20_29_inner_macOut = ($signed(io_mulInput) * $signed(_20_29_inner_activation));
  assign _zz__zz__20_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_29_inner_macOut)) ? 16'h007f : _zz__20_29_inner_macOut_2);
  assign _zz__20_29_inner_macOut_2 = (($signed(_zz__20_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_29_inner_activation;
    end else begin
      io_macOut = _20_29_inner_macOut;
    end
  end

  assign _zz__20_29_inner_macOut = ($signed(_zz__zz__20_29_inner_macOut) + $signed(_zz__zz__20_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_29_inner_activation <= 8'h00;
      _20_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_29_inner_activation <= io_addInput;
      end else begin
        _20_29_inner_macOut <= _zz__20_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_668 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_28_inner_macOut;
  wire       [15:0]   _zz__zz__20_28_inner_macOut_1;
  wire       [15:0]   _zz__20_28_inner_macOut_1;
  wire       [15:0]   _zz__20_28_inner_macOut_2;
  reg        [7:0]    _20_28_inner_activation;
  reg        [7:0]    _20_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_28_inner_macOut;

  assign _zz__zz__20_28_inner_macOut = ($signed(io_mulInput) * $signed(_20_28_inner_activation));
  assign _zz__zz__20_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_28_inner_macOut)) ? 16'h007f : _zz__20_28_inner_macOut_2);
  assign _zz__20_28_inner_macOut_2 = (($signed(_zz__20_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_28_inner_activation;
    end else begin
      io_macOut = _20_28_inner_macOut;
    end
  end

  assign _zz__20_28_inner_macOut = ($signed(_zz__zz__20_28_inner_macOut) + $signed(_zz__zz__20_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_28_inner_activation <= 8'h00;
      _20_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_28_inner_activation <= io_addInput;
      end else begin
        _20_28_inner_macOut <= _zz__20_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_667 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_27_inner_macOut;
  wire       [15:0]   _zz__zz__20_27_inner_macOut_1;
  wire       [15:0]   _zz__20_27_inner_macOut_1;
  wire       [15:0]   _zz__20_27_inner_macOut_2;
  reg        [7:0]    _20_27_inner_activation;
  reg        [7:0]    _20_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_27_inner_macOut;

  assign _zz__zz__20_27_inner_macOut = ($signed(io_mulInput) * $signed(_20_27_inner_activation));
  assign _zz__zz__20_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_27_inner_macOut)) ? 16'h007f : _zz__20_27_inner_macOut_2);
  assign _zz__20_27_inner_macOut_2 = (($signed(_zz__20_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_27_inner_activation;
    end else begin
      io_macOut = _20_27_inner_macOut;
    end
  end

  assign _zz__20_27_inner_macOut = ($signed(_zz__zz__20_27_inner_macOut) + $signed(_zz__zz__20_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_27_inner_activation <= 8'h00;
      _20_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_27_inner_activation <= io_addInput;
      end else begin
        _20_27_inner_macOut <= _zz__20_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_666 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_26_inner_macOut;
  wire       [15:0]   _zz__zz__20_26_inner_macOut_1;
  wire       [15:0]   _zz__20_26_inner_macOut_1;
  wire       [15:0]   _zz__20_26_inner_macOut_2;
  reg        [7:0]    _20_26_inner_activation;
  reg        [7:0]    _20_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_26_inner_macOut;

  assign _zz__zz__20_26_inner_macOut = ($signed(io_mulInput) * $signed(_20_26_inner_activation));
  assign _zz__zz__20_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_26_inner_macOut)) ? 16'h007f : _zz__20_26_inner_macOut_2);
  assign _zz__20_26_inner_macOut_2 = (($signed(_zz__20_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_26_inner_activation;
    end else begin
      io_macOut = _20_26_inner_macOut;
    end
  end

  assign _zz__20_26_inner_macOut = ($signed(_zz__zz__20_26_inner_macOut) + $signed(_zz__zz__20_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_26_inner_activation <= 8'h00;
      _20_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_26_inner_activation <= io_addInput;
      end else begin
        _20_26_inner_macOut <= _zz__20_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_665 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_25_inner_macOut;
  wire       [15:0]   _zz__zz__20_25_inner_macOut_1;
  wire       [15:0]   _zz__20_25_inner_macOut_1;
  wire       [15:0]   _zz__20_25_inner_macOut_2;
  reg        [7:0]    _20_25_inner_activation;
  reg        [7:0]    _20_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_25_inner_macOut;

  assign _zz__zz__20_25_inner_macOut = ($signed(io_mulInput) * $signed(_20_25_inner_activation));
  assign _zz__zz__20_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_25_inner_macOut)) ? 16'h007f : _zz__20_25_inner_macOut_2);
  assign _zz__20_25_inner_macOut_2 = (($signed(_zz__20_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_25_inner_activation;
    end else begin
      io_macOut = _20_25_inner_macOut;
    end
  end

  assign _zz__20_25_inner_macOut = ($signed(_zz__zz__20_25_inner_macOut) + $signed(_zz__zz__20_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_25_inner_activation <= 8'h00;
      _20_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_25_inner_activation <= io_addInput;
      end else begin
        _20_25_inner_macOut <= _zz__20_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_664 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_24_inner_macOut;
  wire       [15:0]   _zz__zz__20_24_inner_macOut_1;
  wire       [15:0]   _zz__20_24_inner_macOut_1;
  wire       [15:0]   _zz__20_24_inner_macOut_2;
  reg        [7:0]    _20_24_inner_activation;
  reg        [7:0]    _20_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_24_inner_macOut;

  assign _zz__zz__20_24_inner_macOut = ($signed(io_mulInput) * $signed(_20_24_inner_activation));
  assign _zz__zz__20_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_24_inner_macOut)) ? 16'h007f : _zz__20_24_inner_macOut_2);
  assign _zz__20_24_inner_macOut_2 = (($signed(_zz__20_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_24_inner_activation;
    end else begin
      io_macOut = _20_24_inner_macOut;
    end
  end

  assign _zz__20_24_inner_macOut = ($signed(_zz__zz__20_24_inner_macOut) + $signed(_zz__zz__20_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_24_inner_activation <= 8'h00;
      _20_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_24_inner_activation <= io_addInput;
      end else begin
        _20_24_inner_macOut <= _zz__20_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_663 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_23_inner_macOut;
  wire       [15:0]   _zz__zz__20_23_inner_macOut_1;
  wire       [15:0]   _zz__20_23_inner_macOut_1;
  wire       [15:0]   _zz__20_23_inner_macOut_2;
  reg        [7:0]    _20_23_inner_activation;
  reg        [7:0]    _20_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_23_inner_macOut;

  assign _zz__zz__20_23_inner_macOut = ($signed(io_mulInput) * $signed(_20_23_inner_activation));
  assign _zz__zz__20_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_23_inner_macOut)) ? 16'h007f : _zz__20_23_inner_macOut_2);
  assign _zz__20_23_inner_macOut_2 = (($signed(_zz__20_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_23_inner_activation;
    end else begin
      io_macOut = _20_23_inner_macOut;
    end
  end

  assign _zz__20_23_inner_macOut = ($signed(_zz__zz__20_23_inner_macOut) + $signed(_zz__zz__20_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_23_inner_activation <= 8'h00;
      _20_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_23_inner_activation <= io_addInput;
      end else begin
        _20_23_inner_macOut <= _zz__20_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_662 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_22_inner_macOut;
  wire       [15:0]   _zz__zz__20_22_inner_macOut_1;
  wire       [15:0]   _zz__20_22_inner_macOut_1;
  wire       [15:0]   _zz__20_22_inner_macOut_2;
  reg        [7:0]    _20_22_inner_activation;
  reg        [7:0]    _20_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_22_inner_macOut;

  assign _zz__zz__20_22_inner_macOut = ($signed(io_mulInput) * $signed(_20_22_inner_activation));
  assign _zz__zz__20_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_22_inner_macOut)) ? 16'h007f : _zz__20_22_inner_macOut_2);
  assign _zz__20_22_inner_macOut_2 = (($signed(_zz__20_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_22_inner_activation;
    end else begin
      io_macOut = _20_22_inner_macOut;
    end
  end

  assign _zz__20_22_inner_macOut = ($signed(_zz__zz__20_22_inner_macOut) + $signed(_zz__zz__20_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_22_inner_activation <= 8'h00;
      _20_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_22_inner_activation <= io_addInput;
      end else begin
        _20_22_inner_macOut <= _zz__20_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_661 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_21_inner_macOut;
  wire       [15:0]   _zz__zz__20_21_inner_macOut_1;
  wire       [15:0]   _zz__20_21_inner_macOut_1;
  wire       [15:0]   _zz__20_21_inner_macOut_2;
  reg        [7:0]    _20_21_inner_activation;
  reg        [7:0]    _20_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_21_inner_macOut;

  assign _zz__zz__20_21_inner_macOut = ($signed(io_mulInput) * $signed(_20_21_inner_activation));
  assign _zz__zz__20_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_21_inner_macOut)) ? 16'h007f : _zz__20_21_inner_macOut_2);
  assign _zz__20_21_inner_macOut_2 = (($signed(_zz__20_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_21_inner_activation;
    end else begin
      io_macOut = _20_21_inner_macOut;
    end
  end

  assign _zz__20_21_inner_macOut = ($signed(_zz__zz__20_21_inner_macOut) + $signed(_zz__zz__20_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_21_inner_activation <= 8'h00;
      _20_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_21_inner_activation <= io_addInput;
      end else begin
        _20_21_inner_macOut <= _zz__20_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_660 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_20_inner_macOut;
  wire       [15:0]   _zz__zz__20_20_inner_macOut_1;
  wire       [15:0]   _zz__20_20_inner_macOut_1;
  wire       [15:0]   _zz__20_20_inner_macOut_2;
  reg        [7:0]    _20_20_inner_activation;
  reg        [7:0]    _20_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_20_inner_macOut;

  assign _zz__zz__20_20_inner_macOut = ($signed(io_mulInput) * $signed(_20_20_inner_activation));
  assign _zz__zz__20_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_20_inner_macOut)) ? 16'h007f : _zz__20_20_inner_macOut_2);
  assign _zz__20_20_inner_macOut_2 = (($signed(_zz__20_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_20_inner_activation;
    end else begin
      io_macOut = _20_20_inner_macOut;
    end
  end

  assign _zz__20_20_inner_macOut = ($signed(_zz__zz__20_20_inner_macOut) + $signed(_zz__zz__20_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_20_inner_activation <= 8'h00;
      _20_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_20_inner_activation <= io_addInput;
      end else begin
        _20_20_inner_macOut <= _zz__20_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_659 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_19_inner_macOut;
  wire       [15:0]   _zz__zz__20_19_inner_macOut_1;
  wire       [15:0]   _zz__20_19_inner_macOut_1;
  wire       [15:0]   _zz__20_19_inner_macOut_2;
  reg        [7:0]    _20_19_inner_activation;
  reg        [7:0]    _20_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_19_inner_macOut;

  assign _zz__zz__20_19_inner_macOut = ($signed(io_mulInput) * $signed(_20_19_inner_activation));
  assign _zz__zz__20_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_19_inner_macOut)) ? 16'h007f : _zz__20_19_inner_macOut_2);
  assign _zz__20_19_inner_macOut_2 = (($signed(_zz__20_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_19_inner_activation;
    end else begin
      io_macOut = _20_19_inner_macOut;
    end
  end

  assign _zz__20_19_inner_macOut = ($signed(_zz__zz__20_19_inner_macOut) + $signed(_zz__zz__20_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_19_inner_activation <= 8'h00;
      _20_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_19_inner_activation <= io_addInput;
      end else begin
        _20_19_inner_macOut <= _zz__20_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_658 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_18_inner_macOut;
  wire       [15:0]   _zz__zz__20_18_inner_macOut_1;
  wire       [15:0]   _zz__20_18_inner_macOut_1;
  wire       [15:0]   _zz__20_18_inner_macOut_2;
  reg        [7:0]    _20_18_inner_activation;
  reg        [7:0]    _20_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_18_inner_macOut;

  assign _zz__zz__20_18_inner_macOut = ($signed(io_mulInput) * $signed(_20_18_inner_activation));
  assign _zz__zz__20_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_18_inner_macOut)) ? 16'h007f : _zz__20_18_inner_macOut_2);
  assign _zz__20_18_inner_macOut_2 = (($signed(_zz__20_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_18_inner_activation;
    end else begin
      io_macOut = _20_18_inner_macOut;
    end
  end

  assign _zz__20_18_inner_macOut = ($signed(_zz__zz__20_18_inner_macOut) + $signed(_zz__zz__20_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_18_inner_activation <= 8'h00;
      _20_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_18_inner_activation <= io_addInput;
      end else begin
        _20_18_inner_macOut <= _zz__20_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_657 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_17_inner_macOut;
  wire       [15:0]   _zz__zz__20_17_inner_macOut_1;
  wire       [15:0]   _zz__20_17_inner_macOut_1;
  wire       [15:0]   _zz__20_17_inner_macOut_2;
  reg        [7:0]    _20_17_inner_activation;
  reg        [7:0]    _20_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_17_inner_macOut;

  assign _zz__zz__20_17_inner_macOut = ($signed(io_mulInput) * $signed(_20_17_inner_activation));
  assign _zz__zz__20_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_17_inner_macOut)) ? 16'h007f : _zz__20_17_inner_macOut_2);
  assign _zz__20_17_inner_macOut_2 = (($signed(_zz__20_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_17_inner_activation;
    end else begin
      io_macOut = _20_17_inner_macOut;
    end
  end

  assign _zz__20_17_inner_macOut = ($signed(_zz__zz__20_17_inner_macOut) + $signed(_zz__zz__20_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_17_inner_activation <= 8'h00;
      _20_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_17_inner_activation <= io_addInput;
      end else begin
        _20_17_inner_macOut <= _zz__20_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_656 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_16_inner_macOut;
  wire       [15:0]   _zz__zz__20_16_inner_macOut_1;
  wire       [15:0]   _zz__20_16_inner_macOut_1;
  wire       [15:0]   _zz__20_16_inner_macOut_2;
  reg        [7:0]    _20_16_inner_activation;
  reg        [7:0]    _20_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_16_inner_macOut;

  assign _zz__zz__20_16_inner_macOut = ($signed(io_mulInput) * $signed(_20_16_inner_activation));
  assign _zz__zz__20_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_16_inner_macOut)) ? 16'h007f : _zz__20_16_inner_macOut_2);
  assign _zz__20_16_inner_macOut_2 = (($signed(_zz__20_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_16_inner_activation;
    end else begin
      io_macOut = _20_16_inner_macOut;
    end
  end

  assign _zz__20_16_inner_macOut = ($signed(_zz__zz__20_16_inner_macOut) + $signed(_zz__zz__20_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_16_inner_activation <= 8'h00;
      _20_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_16_inner_activation <= io_addInput;
      end else begin
        _20_16_inner_macOut <= _zz__20_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_655 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_15_inner_macOut;
  wire       [15:0]   _zz__zz__20_15_inner_macOut_1;
  wire       [15:0]   _zz__20_15_inner_macOut_1;
  wire       [15:0]   _zz__20_15_inner_macOut_2;
  reg        [7:0]    _20_15_inner_activation;
  reg        [7:0]    _20_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_15_inner_macOut;

  assign _zz__zz__20_15_inner_macOut = ($signed(io_mulInput) * $signed(_20_15_inner_activation));
  assign _zz__zz__20_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_15_inner_macOut)) ? 16'h007f : _zz__20_15_inner_macOut_2);
  assign _zz__20_15_inner_macOut_2 = (($signed(_zz__20_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_15_inner_activation;
    end else begin
      io_macOut = _20_15_inner_macOut;
    end
  end

  assign _zz__20_15_inner_macOut = ($signed(_zz__zz__20_15_inner_macOut) + $signed(_zz__zz__20_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_15_inner_activation <= 8'h00;
      _20_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_15_inner_activation <= io_addInput;
      end else begin
        _20_15_inner_macOut <= _zz__20_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_654 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_14_inner_macOut;
  wire       [15:0]   _zz__zz__20_14_inner_macOut_1;
  wire       [15:0]   _zz__20_14_inner_macOut_1;
  wire       [15:0]   _zz__20_14_inner_macOut_2;
  reg        [7:0]    _20_14_inner_activation;
  reg        [7:0]    _20_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_14_inner_macOut;

  assign _zz__zz__20_14_inner_macOut = ($signed(io_mulInput) * $signed(_20_14_inner_activation));
  assign _zz__zz__20_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_14_inner_macOut)) ? 16'h007f : _zz__20_14_inner_macOut_2);
  assign _zz__20_14_inner_macOut_2 = (($signed(_zz__20_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_14_inner_activation;
    end else begin
      io_macOut = _20_14_inner_macOut;
    end
  end

  assign _zz__20_14_inner_macOut = ($signed(_zz__zz__20_14_inner_macOut) + $signed(_zz__zz__20_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_14_inner_activation <= 8'h00;
      _20_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_14_inner_activation <= io_addInput;
      end else begin
        _20_14_inner_macOut <= _zz__20_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_653 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_13_inner_macOut;
  wire       [15:0]   _zz__zz__20_13_inner_macOut_1;
  wire       [15:0]   _zz__20_13_inner_macOut_1;
  wire       [15:0]   _zz__20_13_inner_macOut_2;
  reg        [7:0]    _20_13_inner_activation;
  reg        [7:0]    _20_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_13_inner_macOut;

  assign _zz__zz__20_13_inner_macOut = ($signed(io_mulInput) * $signed(_20_13_inner_activation));
  assign _zz__zz__20_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_13_inner_macOut)) ? 16'h007f : _zz__20_13_inner_macOut_2);
  assign _zz__20_13_inner_macOut_2 = (($signed(_zz__20_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_13_inner_activation;
    end else begin
      io_macOut = _20_13_inner_macOut;
    end
  end

  assign _zz__20_13_inner_macOut = ($signed(_zz__zz__20_13_inner_macOut) + $signed(_zz__zz__20_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_13_inner_activation <= 8'h00;
      _20_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_13_inner_activation <= io_addInput;
      end else begin
        _20_13_inner_macOut <= _zz__20_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_652 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_12_inner_macOut;
  wire       [15:0]   _zz__zz__20_12_inner_macOut_1;
  wire       [15:0]   _zz__20_12_inner_macOut_1;
  wire       [15:0]   _zz__20_12_inner_macOut_2;
  reg        [7:0]    _20_12_inner_activation;
  reg        [7:0]    _20_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_12_inner_macOut;

  assign _zz__zz__20_12_inner_macOut = ($signed(io_mulInput) * $signed(_20_12_inner_activation));
  assign _zz__zz__20_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_12_inner_macOut)) ? 16'h007f : _zz__20_12_inner_macOut_2);
  assign _zz__20_12_inner_macOut_2 = (($signed(_zz__20_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_12_inner_activation;
    end else begin
      io_macOut = _20_12_inner_macOut;
    end
  end

  assign _zz__20_12_inner_macOut = ($signed(_zz__zz__20_12_inner_macOut) + $signed(_zz__zz__20_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_12_inner_activation <= 8'h00;
      _20_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_12_inner_activation <= io_addInput;
      end else begin
        _20_12_inner_macOut <= _zz__20_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_651 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_11_inner_macOut;
  wire       [15:0]   _zz__zz__20_11_inner_macOut_1;
  wire       [15:0]   _zz__20_11_inner_macOut_1;
  wire       [15:0]   _zz__20_11_inner_macOut_2;
  reg        [7:0]    _20_11_inner_activation;
  reg        [7:0]    _20_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_11_inner_macOut;

  assign _zz__zz__20_11_inner_macOut = ($signed(io_mulInput) * $signed(_20_11_inner_activation));
  assign _zz__zz__20_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_11_inner_macOut)) ? 16'h007f : _zz__20_11_inner_macOut_2);
  assign _zz__20_11_inner_macOut_2 = (($signed(_zz__20_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_11_inner_activation;
    end else begin
      io_macOut = _20_11_inner_macOut;
    end
  end

  assign _zz__20_11_inner_macOut = ($signed(_zz__zz__20_11_inner_macOut) + $signed(_zz__zz__20_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_11_inner_activation <= 8'h00;
      _20_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_11_inner_activation <= io_addInput;
      end else begin
        _20_11_inner_macOut <= _zz__20_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_650 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_10_inner_macOut;
  wire       [15:0]   _zz__zz__20_10_inner_macOut_1;
  wire       [15:0]   _zz__20_10_inner_macOut_1;
  wire       [15:0]   _zz__20_10_inner_macOut_2;
  reg        [7:0]    _20_10_inner_activation;
  reg        [7:0]    _20_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_10_inner_macOut;

  assign _zz__zz__20_10_inner_macOut = ($signed(io_mulInput) * $signed(_20_10_inner_activation));
  assign _zz__zz__20_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_10_inner_macOut)) ? 16'h007f : _zz__20_10_inner_macOut_2);
  assign _zz__20_10_inner_macOut_2 = (($signed(_zz__20_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_10_inner_activation;
    end else begin
      io_macOut = _20_10_inner_macOut;
    end
  end

  assign _zz__20_10_inner_macOut = ($signed(_zz__zz__20_10_inner_macOut) + $signed(_zz__zz__20_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_10_inner_activation <= 8'h00;
      _20_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_10_inner_activation <= io_addInput;
      end else begin
        _20_10_inner_macOut <= _zz__20_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_649 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_9_inner_macOut;
  wire       [15:0]   _zz__zz__20_9_inner_macOut_1;
  wire       [15:0]   _zz__20_9_inner_macOut_1;
  wire       [15:0]   _zz__20_9_inner_macOut_2;
  reg        [7:0]    _20_9_inner_activation;
  reg        [7:0]    _20_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_9_inner_macOut;

  assign _zz__zz__20_9_inner_macOut = ($signed(io_mulInput) * $signed(_20_9_inner_activation));
  assign _zz__zz__20_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_9_inner_macOut)) ? 16'h007f : _zz__20_9_inner_macOut_2);
  assign _zz__20_9_inner_macOut_2 = (($signed(_zz__20_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_9_inner_activation;
    end else begin
      io_macOut = _20_9_inner_macOut;
    end
  end

  assign _zz__20_9_inner_macOut = ($signed(_zz__zz__20_9_inner_macOut) + $signed(_zz__zz__20_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_9_inner_activation <= 8'h00;
      _20_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_9_inner_activation <= io_addInput;
      end else begin
        _20_9_inner_macOut <= _zz__20_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_648 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_8_inner_macOut;
  wire       [15:0]   _zz__zz__20_8_inner_macOut_1;
  wire       [15:0]   _zz__20_8_inner_macOut_1;
  wire       [15:0]   _zz__20_8_inner_macOut_2;
  reg        [7:0]    _20_8_inner_activation;
  reg        [7:0]    _20_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_8_inner_macOut;

  assign _zz__zz__20_8_inner_macOut = ($signed(io_mulInput) * $signed(_20_8_inner_activation));
  assign _zz__zz__20_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_8_inner_macOut)) ? 16'h007f : _zz__20_8_inner_macOut_2);
  assign _zz__20_8_inner_macOut_2 = (($signed(_zz__20_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_8_inner_activation;
    end else begin
      io_macOut = _20_8_inner_macOut;
    end
  end

  assign _zz__20_8_inner_macOut = ($signed(_zz__zz__20_8_inner_macOut) + $signed(_zz__zz__20_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_8_inner_activation <= 8'h00;
      _20_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_8_inner_activation <= io_addInput;
      end else begin
        _20_8_inner_macOut <= _zz__20_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_647 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_7_inner_macOut;
  wire       [15:0]   _zz__zz__20_7_inner_macOut_1;
  wire       [15:0]   _zz__20_7_inner_macOut_1;
  wire       [15:0]   _zz__20_7_inner_macOut_2;
  reg        [7:0]    _20_7_inner_activation;
  reg        [7:0]    _20_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_7_inner_macOut;

  assign _zz__zz__20_7_inner_macOut = ($signed(io_mulInput) * $signed(_20_7_inner_activation));
  assign _zz__zz__20_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_7_inner_macOut)) ? 16'h007f : _zz__20_7_inner_macOut_2);
  assign _zz__20_7_inner_macOut_2 = (($signed(_zz__20_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_7_inner_activation;
    end else begin
      io_macOut = _20_7_inner_macOut;
    end
  end

  assign _zz__20_7_inner_macOut = ($signed(_zz__zz__20_7_inner_macOut) + $signed(_zz__zz__20_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_7_inner_activation <= 8'h00;
      _20_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_7_inner_activation <= io_addInput;
      end else begin
        _20_7_inner_macOut <= _zz__20_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_646 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_6_inner_macOut;
  wire       [15:0]   _zz__zz__20_6_inner_macOut_1;
  wire       [15:0]   _zz__20_6_inner_macOut_1;
  wire       [15:0]   _zz__20_6_inner_macOut_2;
  reg        [7:0]    _20_6_inner_activation;
  reg        [7:0]    _20_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_6_inner_macOut;

  assign _zz__zz__20_6_inner_macOut = ($signed(io_mulInput) * $signed(_20_6_inner_activation));
  assign _zz__zz__20_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_6_inner_macOut)) ? 16'h007f : _zz__20_6_inner_macOut_2);
  assign _zz__20_6_inner_macOut_2 = (($signed(_zz__20_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_6_inner_activation;
    end else begin
      io_macOut = _20_6_inner_macOut;
    end
  end

  assign _zz__20_6_inner_macOut = ($signed(_zz__zz__20_6_inner_macOut) + $signed(_zz__zz__20_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_6_inner_activation <= 8'h00;
      _20_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_6_inner_activation <= io_addInput;
      end else begin
        _20_6_inner_macOut <= _zz__20_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_645 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_5_inner_macOut;
  wire       [15:0]   _zz__zz__20_5_inner_macOut_1;
  wire       [15:0]   _zz__20_5_inner_macOut_1;
  wire       [15:0]   _zz__20_5_inner_macOut_2;
  reg        [7:0]    _20_5_inner_activation;
  reg        [7:0]    _20_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_5_inner_macOut;

  assign _zz__zz__20_5_inner_macOut = ($signed(io_mulInput) * $signed(_20_5_inner_activation));
  assign _zz__zz__20_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_5_inner_macOut)) ? 16'h007f : _zz__20_5_inner_macOut_2);
  assign _zz__20_5_inner_macOut_2 = (($signed(_zz__20_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_5_inner_activation;
    end else begin
      io_macOut = _20_5_inner_macOut;
    end
  end

  assign _zz__20_5_inner_macOut = ($signed(_zz__zz__20_5_inner_macOut) + $signed(_zz__zz__20_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_5_inner_activation <= 8'h00;
      _20_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_5_inner_activation <= io_addInput;
      end else begin
        _20_5_inner_macOut <= _zz__20_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_644 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_4_inner_macOut;
  wire       [15:0]   _zz__zz__20_4_inner_macOut_1;
  wire       [15:0]   _zz__20_4_inner_macOut_1;
  wire       [15:0]   _zz__20_4_inner_macOut_2;
  reg        [7:0]    _20_4_inner_activation;
  reg        [7:0]    _20_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_4_inner_macOut;

  assign _zz__zz__20_4_inner_macOut = ($signed(io_mulInput) * $signed(_20_4_inner_activation));
  assign _zz__zz__20_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_4_inner_macOut)) ? 16'h007f : _zz__20_4_inner_macOut_2);
  assign _zz__20_4_inner_macOut_2 = (($signed(_zz__20_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_4_inner_activation;
    end else begin
      io_macOut = _20_4_inner_macOut;
    end
  end

  assign _zz__20_4_inner_macOut = ($signed(_zz__zz__20_4_inner_macOut) + $signed(_zz__zz__20_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_4_inner_activation <= 8'h00;
      _20_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_4_inner_activation <= io_addInput;
      end else begin
        _20_4_inner_macOut <= _zz__20_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_643 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_3_inner_macOut;
  wire       [15:0]   _zz__zz__20_3_inner_macOut_1;
  wire       [15:0]   _zz__20_3_inner_macOut_1;
  wire       [15:0]   _zz__20_3_inner_macOut_2;
  reg        [7:0]    _20_3_inner_activation;
  reg        [7:0]    _20_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_3_inner_macOut;

  assign _zz__zz__20_3_inner_macOut = ($signed(io_mulInput) * $signed(_20_3_inner_activation));
  assign _zz__zz__20_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_3_inner_macOut)) ? 16'h007f : _zz__20_3_inner_macOut_2);
  assign _zz__20_3_inner_macOut_2 = (($signed(_zz__20_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_3_inner_activation;
    end else begin
      io_macOut = _20_3_inner_macOut;
    end
  end

  assign _zz__20_3_inner_macOut = ($signed(_zz__zz__20_3_inner_macOut) + $signed(_zz__zz__20_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_3_inner_activation <= 8'h00;
      _20_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_3_inner_activation <= io_addInput;
      end else begin
        _20_3_inner_macOut <= _zz__20_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_642 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_2_inner_macOut;
  wire       [15:0]   _zz__zz__20_2_inner_macOut_1;
  wire       [15:0]   _zz__20_2_inner_macOut_1;
  wire       [15:0]   _zz__20_2_inner_macOut_2;
  reg        [7:0]    _20_2_inner_activation;
  reg        [7:0]    _20_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_2_inner_macOut;

  assign _zz__zz__20_2_inner_macOut = ($signed(io_mulInput) * $signed(_20_2_inner_activation));
  assign _zz__zz__20_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_2_inner_macOut)) ? 16'h007f : _zz__20_2_inner_macOut_2);
  assign _zz__20_2_inner_macOut_2 = (($signed(_zz__20_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_2_inner_activation;
    end else begin
      io_macOut = _20_2_inner_macOut;
    end
  end

  assign _zz__20_2_inner_macOut = ($signed(_zz__zz__20_2_inner_macOut) + $signed(_zz__zz__20_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_2_inner_activation <= 8'h00;
      _20_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_2_inner_activation <= io_addInput;
      end else begin
        _20_2_inner_macOut <= _zz__20_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_641 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_1_inner_macOut;
  wire       [15:0]   _zz__zz__20_1_inner_macOut_1;
  wire       [15:0]   _zz__20_1_inner_macOut_1;
  wire       [15:0]   _zz__20_1_inner_macOut_2;
  reg        [7:0]    _20_1_inner_activation;
  reg        [7:0]    _20_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_1_inner_macOut;

  assign _zz__zz__20_1_inner_macOut = ($signed(io_mulInput) * $signed(_20_1_inner_activation));
  assign _zz__zz__20_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_1_inner_macOut)) ? 16'h007f : _zz__20_1_inner_macOut_2);
  assign _zz__20_1_inner_macOut_2 = (($signed(_zz__20_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_1_inner_activation;
    end else begin
      io_macOut = _20_1_inner_macOut;
    end
  end

  assign _zz__20_1_inner_macOut = ($signed(_zz__zz__20_1_inner_macOut) + $signed(_zz__zz__20_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_1_inner_activation <= 8'h00;
      _20_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_1_inner_activation <= io_addInput;
      end else begin
        _20_1_inner_macOut <= _zz__20_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_640 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__20_0_inner_macOut;
  wire       [15:0]   _zz__zz__20_0_inner_macOut_1;
  wire       [15:0]   _zz__20_0_inner_macOut_1;
  wire       [15:0]   _zz__20_0_inner_macOut_2;
  reg        [7:0]    _20_0_inner_activation;
  reg        [7:0]    _20_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__20_0_inner_macOut;

  assign _zz__zz__20_0_inner_macOut = ($signed(io_mulInput) * $signed(_20_0_inner_activation));
  assign _zz__zz__20_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__20_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__20_0_inner_macOut)) ? 16'h007f : _zz__20_0_inner_macOut_2);
  assign _zz__20_0_inner_macOut_2 = (($signed(_zz__20_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__20_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _20_0_inner_activation;
    end else begin
      io_macOut = _20_0_inner_macOut;
    end
  end

  assign _zz__20_0_inner_macOut = ($signed(_zz__zz__20_0_inner_macOut) + $signed(_zz__zz__20_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _20_0_inner_activation <= 8'h00;
      _20_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _20_0_inner_activation <= io_addInput;
      end else begin
        _20_0_inner_macOut <= _zz__20_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_639 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_31_inner_macOut;
  wire       [15:0]   _zz__zz__19_31_inner_macOut_1;
  wire       [15:0]   _zz__19_31_inner_macOut_1;
  wire       [15:0]   _zz__19_31_inner_macOut_2;
  reg        [7:0]    _19_31_inner_activation;
  reg        [7:0]    _19_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_31_inner_macOut;

  assign _zz__zz__19_31_inner_macOut = ($signed(io_mulInput) * $signed(_19_31_inner_activation));
  assign _zz__zz__19_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_31_inner_macOut)) ? 16'h007f : _zz__19_31_inner_macOut_2);
  assign _zz__19_31_inner_macOut_2 = (($signed(_zz__19_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_31_inner_activation;
    end else begin
      io_macOut = _19_31_inner_macOut;
    end
  end

  assign _zz__19_31_inner_macOut = ($signed(_zz__zz__19_31_inner_macOut) + $signed(_zz__zz__19_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_31_inner_activation <= 8'h00;
      _19_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_31_inner_activation <= io_addInput;
      end else begin
        _19_31_inner_macOut <= _zz__19_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_638 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_30_inner_macOut;
  wire       [15:0]   _zz__zz__19_30_inner_macOut_1;
  wire       [15:0]   _zz__19_30_inner_macOut_1;
  wire       [15:0]   _zz__19_30_inner_macOut_2;
  reg        [7:0]    _19_30_inner_activation;
  reg        [7:0]    _19_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_30_inner_macOut;

  assign _zz__zz__19_30_inner_macOut = ($signed(io_mulInput) * $signed(_19_30_inner_activation));
  assign _zz__zz__19_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_30_inner_macOut)) ? 16'h007f : _zz__19_30_inner_macOut_2);
  assign _zz__19_30_inner_macOut_2 = (($signed(_zz__19_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_30_inner_activation;
    end else begin
      io_macOut = _19_30_inner_macOut;
    end
  end

  assign _zz__19_30_inner_macOut = ($signed(_zz__zz__19_30_inner_macOut) + $signed(_zz__zz__19_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_30_inner_activation <= 8'h00;
      _19_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_30_inner_activation <= io_addInput;
      end else begin
        _19_30_inner_macOut <= _zz__19_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_637 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_29_inner_macOut;
  wire       [15:0]   _zz__zz__19_29_inner_macOut_1;
  wire       [15:0]   _zz__19_29_inner_macOut_1;
  wire       [15:0]   _zz__19_29_inner_macOut_2;
  reg        [7:0]    _19_29_inner_activation;
  reg        [7:0]    _19_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_29_inner_macOut;

  assign _zz__zz__19_29_inner_macOut = ($signed(io_mulInput) * $signed(_19_29_inner_activation));
  assign _zz__zz__19_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_29_inner_macOut)) ? 16'h007f : _zz__19_29_inner_macOut_2);
  assign _zz__19_29_inner_macOut_2 = (($signed(_zz__19_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_29_inner_activation;
    end else begin
      io_macOut = _19_29_inner_macOut;
    end
  end

  assign _zz__19_29_inner_macOut = ($signed(_zz__zz__19_29_inner_macOut) + $signed(_zz__zz__19_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_29_inner_activation <= 8'h00;
      _19_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_29_inner_activation <= io_addInput;
      end else begin
        _19_29_inner_macOut <= _zz__19_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_636 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_28_inner_macOut;
  wire       [15:0]   _zz__zz__19_28_inner_macOut_1;
  wire       [15:0]   _zz__19_28_inner_macOut_1;
  wire       [15:0]   _zz__19_28_inner_macOut_2;
  reg        [7:0]    _19_28_inner_activation;
  reg        [7:0]    _19_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_28_inner_macOut;

  assign _zz__zz__19_28_inner_macOut = ($signed(io_mulInput) * $signed(_19_28_inner_activation));
  assign _zz__zz__19_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_28_inner_macOut)) ? 16'h007f : _zz__19_28_inner_macOut_2);
  assign _zz__19_28_inner_macOut_2 = (($signed(_zz__19_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_28_inner_activation;
    end else begin
      io_macOut = _19_28_inner_macOut;
    end
  end

  assign _zz__19_28_inner_macOut = ($signed(_zz__zz__19_28_inner_macOut) + $signed(_zz__zz__19_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_28_inner_activation <= 8'h00;
      _19_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_28_inner_activation <= io_addInput;
      end else begin
        _19_28_inner_macOut <= _zz__19_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_635 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_27_inner_macOut;
  wire       [15:0]   _zz__zz__19_27_inner_macOut_1;
  wire       [15:0]   _zz__19_27_inner_macOut_1;
  wire       [15:0]   _zz__19_27_inner_macOut_2;
  reg        [7:0]    _19_27_inner_activation;
  reg        [7:0]    _19_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_27_inner_macOut;

  assign _zz__zz__19_27_inner_macOut = ($signed(io_mulInput) * $signed(_19_27_inner_activation));
  assign _zz__zz__19_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_27_inner_macOut)) ? 16'h007f : _zz__19_27_inner_macOut_2);
  assign _zz__19_27_inner_macOut_2 = (($signed(_zz__19_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_27_inner_activation;
    end else begin
      io_macOut = _19_27_inner_macOut;
    end
  end

  assign _zz__19_27_inner_macOut = ($signed(_zz__zz__19_27_inner_macOut) + $signed(_zz__zz__19_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_27_inner_activation <= 8'h00;
      _19_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_27_inner_activation <= io_addInput;
      end else begin
        _19_27_inner_macOut <= _zz__19_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_634 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_26_inner_macOut;
  wire       [15:0]   _zz__zz__19_26_inner_macOut_1;
  wire       [15:0]   _zz__19_26_inner_macOut_1;
  wire       [15:0]   _zz__19_26_inner_macOut_2;
  reg        [7:0]    _19_26_inner_activation;
  reg        [7:0]    _19_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_26_inner_macOut;

  assign _zz__zz__19_26_inner_macOut = ($signed(io_mulInput) * $signed(_19_26_inner_activation));
  assign _zz__zz__19_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_26_inner_macOut)) ? 16'h007f : _zz__19_26_inner_macOut_2);
  assign _zz__19_26_inner_macOut_2 = (($signed(_zz__19_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_26_inner_activation;
    end else begin
      io_macOut = _19_26_inner_macOut;
    end
  end

  assign _zz__19_26_inner_macOut = ($signed(_zz__zz__19_26_inner_macOut) + $signed(_zz__zz__19_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_26_inner_activation <= 8'h00;
      _19_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_26_inner_activation <= io_addInput;
      end else begin
        _19_26_inner_macOut <= _zz__19_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_633 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_25_inner_macOut;
  wire       [15:0]   _zz__zz__19_25_inner_macOut_1;
  wire       [15:0]   _zz__19_25_inner_macOut_1;
  wire       [15:0]   _zz__19_25_inner_macOut_2;
  reg        [7:0]    _19_25_inner_activation;
  reg        [7:0]    _19_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_25_inner_macOut;

  assign _zz__zz__19_25_inner_macOut = ($signed(io_mulInput) * $signed(_19_25_inner_activation));
  assign _zz__zz__19_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_25_inner_macOut)) ? 16'h007f : _zz__19_25_inner_macOut_2);
  assign _zz__19_25_inner_macOut_2 = (($signed(_zz__19_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_25_inner_activation;
    end else begin
      io_macOut = _19_25_inner_macOut;
    end
  end

  assign _zz__19_25_inner_macOut = ($signed(_zz__zz__19_25_inner_macOut) + $signed(_zz__zz__19_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_25_inner_activation <= 8'h00;
      _19_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_25_inner_activation <= io_addInput;
      end else begin
        _19_25_inner_macOut <= _zz__19_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_632 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_24_inner_macOut;
  wire       [15:0]   _zz__zz__19_24_inner_macOut_1;
  wire       [15:0]   _zz__19_24_inner_macOut_1;
  wire       [15:0]   _zz__19_24_inner_macOut_2;
  reg        [7:0]    _19_24_inner_activation;
  reg        [7:0]    _19_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_24_inner_macOut;

  assign _zz__zz__19_24_inner_macOut = ($signed(io_mulInput) * $signed(_19_24_inner_activation));
  assign _zz__zz__19_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_24_inner_macOut)) ? 16'h007f : _zz__19_24_inner_macOut_2);
  assign _zz__19_24_inner_macOut_2 = (($signed(_zz__19_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_24_inner_activation;
    end else begin
      io_macOut = _19_24_inner_macOut;
    end
  end

  assign _zz__19_24_inner_macOut = ($signed(_zz__zz__19_24_inner_macOut) + $signed(_zz__zz__19_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_24_inner_activation <= 8'h00;
      _19_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_24_inner_activation <= io_addInput;
      end else begin
        _19_24_inner_macOut <= _zz__19_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_631 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_23_inner_macOut;
  wire       [15:0]   _zz__zz__19_23_inner_macOut_1;
  wire       [15:0]   _zz__19_23_inner_macOut_1;
  wire       [15:0]   _zz__19_23_inner_macOut_2;
  reg        [7:0]    _19_23_inner_activation;
  reg        [7:0]    _19_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_23_inner_macOut;

  assign _zz__zz__19_23_inner_macOut = ($signed(io_mulInput) * $signed(_19_23_inner_activation));
  assign _zz__zz__19_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_23_inner_macOut)) ? 16'h007f : _zz__19_23_inner_macOut_2);
  assign _zz__19_23_inner_macOut_2 = (($signed(_zz__19_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_23_inner_activation;
    end else begin
      io_macOut = _19_23_inner_macOut;
    end
  end

  assign _zz__19_23_inner_macOut = ($signed(_zz__zz__19_23_inner_macOut) + $signed(_zz__zz__19_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_23_inner_activation <= 8'h00;
      _19_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_23_inner_activation <= io_addInput;
      end else begin
        _19_23_inner_macOut <= _zz__19_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_630 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_22_inner_macOut;
  wire       [15:0]   _zz__zz__19_22_inner_macOut_1;
  wire       [15:0]   _zz__19_22_inner_macOut_1;
  wire       [15:0]   _zz__19_22_inner_macOut_2;
  reg        [7:0]    _19_22_inner_activation;
  reg        [7:0]    _19_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_22_inner_macOut;

  assign _zz__zz__19_22_inner_macOut = ($signed(io_mulInput) * $signed(_19_22_inner_activation));
  assign _zz__zz__19_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_22_inner_macOut)) ? 16'h007f : _zz__19_22_inner_macOut_2);
  assign _zz__19_22_inner_macOut_2 = (($signed(_zz__19_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_22_inner_activation;
    end else begin
      io_macOut = _19_22_inner_macOut;
    end
  end

  assign _zz__19_22_inner_macOut = ($signed(_zz__zz__19_22_inner_macOut) + $signed(_zz__zz__19_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_22_inner_activation <= 8'h00;
      _19_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_22_inner_activation <= io_addInput;
      end else begin
        _19_22_inner_macOut <= _zz__19_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_629 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_21_inner_macOut;
  wire       [15:0]   _zz__zz__19_21_inner_macOut_1;
  wire       [15:0]   _zz__19_21_inner_macOut_1;
  wire       [15:0]   _zz__19_21_inner_macOut_2;
  reg        [7:0]    _19_21_inner_activation;
  reg        [7:0]    _19_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_21_inner_macOut;

  assign _zz__zz__19_21_inner_macOut = ($signed(io_mulInput) * $signed(_19_21_inner_activation));
  assign _zz__zz__19_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_21_inner_macOut)) ? 16'h007f : _zz__19_21_inner_macOut_2);
  assign _zz__19_21_inner_macOut_2 = (($signed(_zz__19_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_21_inner_activation;
    end else begin
      io_macOut = _19_21_inner_macOut;
    end
  end

  assign _zz__19_21_inner_macOut = ($signed(_zz__zz__19_21_inner_macOut) + $signed(_zz__zz__19_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_21_inner_activation <= 8'h00;
      _19_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_21_inner_activation <= io_addInput;
      end else begin
        _19_21_inner_macOut <= _zz__19_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_628 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_20_inner_macOut;
  wire       [15:0]   _zz__zz__19_20_inner_macOut_1;
  wire       [15:0]   _zz__19_20_inner_macOut_1;
  wire       [15:0]   _zz__19_20_inner_macOut_2;
  reg        [7:0]    _19_20_inner_activation;
  reg        [7:0]    _19_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_20_inner_macOut;

  assign _zz__zz__19_20_inner_macOut = ($signed(io_mulInput) * $signed(_19_20_inner_activation));
  assign _zz__zz__19_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_20_inner_macOut)) ? 16'h007f : _zz__19_20_inner_macOut_2);
  assign _zz__19_20_inner_macOut_2 = (($signed(_zz__19_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_20_inner_activation;
    end else begin
      io_macOut = _19_20_inner_macOut;
    end
  end

  assign _zz__19_20_inner_macOut = ($signed(_zz__zz__19_20_inner_macOut) + $signed(_zz__zz__19_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_20_inner_activation <= 8'h00;
      _19_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_20_inner_activation <= io_addInput;
      end else begin
        _19_20_inner_macOut <= _zz__19_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_627 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_19_inner_macOut;
  wire       [15:0]   _zz__zz__19_19_inner_macOut_1;
  wire       [15:0]   _zz__19_19_inner_macOut_1;
  wire       [15:0]   _zz__19_19_inner_macOut_2;
  reg        [7:0]    _19_19_inner_activation;
  reg        [7:0]    _19_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_19_inner_macOut;

  assign _zz__zz__19_19_inner_macOut = ($signed(io_mulInput) * $signed(_19_19_inner_activation));
  assign _zz__zz__19_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_19_inner_macOut)) ? 16'h007f : _zz__19_19_inner_macOut_2);
  assign _zz__19_19_inner_macOut_2 = (($signed(_zz__19_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_19_inner_activation;
    end else begin
      io_macOut = _19_19_inner_macOut;
    end
  end

  assign _zz__19_19_inner_macOut = ($signed(_zz__zz__19_19_inner_macOut) + $signed(_zz__zz__19_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_19_inner_activation <= 8'h00;
      _19_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_19_inner_activation <= io_addInput;
      end else begin
        _19_19_inner_macOut <= _zz__19_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_626 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_18_inner_macOut;
  wire       [15:0]   _zz__zz__19_18_inner_macOut_1;
  wire       [15:0]   _zz__19_18_inner_macOut_1;
  wire       [15:0]   _zz__19_18_inner_macOut_2;
  reg        [7:0]    _19_18_inner_activation;
  reg        [7:0]    _19_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_18_inner_macOut;

  assign _zz__zz__19_18_inner_macOut = ($signed(io_mulInput) * $signed(_19_18_inner_activation));
  assign _zz__zz__19_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_18_inner_macOut)) ? 16'h007f : _zz__19_18_inner_macOut_2);
  assign _zz__19_18_inner_macOut_2 = (($signed(_zz__19_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_18_inner_activation;
    end else begin
      io_macOut = _19_18_inner_macOut;
    end
  end

  assign _zz__19_18_inner_macOut = ($signed(_zz__zz__19_18_inner_macOut) + $signed(_zz__zz__19_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_18_inner_activation <= 8'h00;
      _19_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_18_inner_activation <= io_addInput;
      end else begin
        _19_18_inner_macOut <= _zz__19_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_625 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_17_inner_macOut;
  wire       [15:0]   _zz__zz__19_17_inner_macOut_1;
  wire       [15:0]   _zz__19_17_inner_macOut_1;
  wire       [15:0]   _zz__19_17_inner_macOut_2;
  reg        [7:0]    _19_17_inner_activation;
  reg        [7:0]    _19_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_17_inner_macOut;

  assign _zz__zz__19_17_inner_macOut = ($signed(io_mulInput) * $signed(_19_17_inner_activation));
  assign _zz__zz__19_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_17_inner_macOut)) ? 16'h007f : _zz__19_17_inner_macOut_2);
  assign _zz__19_17_inner_macOut_2 = (($signed(_zz__19_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_17_inner_activation;
    end else begin
      io_macOut = _19_17_inner_macOut;
    end
  end

  assign _zz__19_17_inner_macOut = ($signed(_zz__zz__19_17_inner_macOut) + $signed(_zz__zz__19_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_17_inner_activation <= 8'h00;
      _19_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_17_inner_activation <= io_addInput;
      end else begin
        _19_17_inner_macOut <= _zz__19_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_624 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_16_inner_macOut;
  wire       [15:0]   _zz__zz__19_16_inner_macOut_1;
  wire       [15:0]   _zz__19_16_inner_macOut_1;
  wire       [15:0]   _zz__19_16_inner_macOut_2;
  reg        [7:0]    _19_16_inner_activation;
  reg        [7:0]    _19_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_16_inner_macOut;

  assign _zz__zz__19_16_inner_macOut = ($signed(io_mulInput) * $signed(_19_16_inner_activation));
  assign _zz__zz__19_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_16_inner_macOut)) ? 16'h007f : _zz__19_16_inner_macOut_2);
  assign _zz__19_16_inner_macOut_2 = (($signed(_zz__19_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_16_inner_activation;
    end else begin
      io_macOut = _19_16_inner_macOut;
    end
  end

  assign _zz__19_16_inner_macOut = ($signed(_zz__zz__19_16_inner_macOut) + $signed(_zz__zz__19_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_16_inner_activation <= 8'h00;
      _19_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_16_inner_activation <= io_addInput;
      end else begin
        _19_16_inner_macOut <= _zz__19_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_623 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_15_inner_macOut;
  wire       [15:0]   _zz__zz__19_15_inner_macOut_1;
  wire       [15:0]   _zz__19_15_inner_macOut_1;
  wire       [15:0]   _zz__19_15_inner_macOut_2;
  reg        [7:0]    _19_15_inner_activation;
  reg        [7:0]    _19_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_15_inner_macOut;

  assign _zz__zz__19_15_inner_macOut = ($signed(io_mulInput) * $signed(_19_15_inner_activation));
  assign _zz__zz__19_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_15_inner_macOut)) ? 16'h007f : _zz__19_15_inner_macOut_2);
  assign _zz__19_15_inner_macOut_2 = (($signed(_zz__19_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_15_inner_activation;
    end else begin
      io_macOut = _19_15_inner_macOut;
    end
  end

  assign _zz__19_15_inner_macOut = ($signed(_zz__zz__19_15_inner_macOut) + $signed(_zz__zz__19_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_15_inner_activation <= 8'h00;
      _19_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_15_inner_activation <= io_addInput;
      end else begin
        _19_15_inner_macOut <= _zz__19_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_622 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_14_inner_macOut;
  wire       [15:0]   _zz__zz__19_14_inner_macOut_1;
  wire       [15:0]   _zz__19_14_inner_macOut_1;
  wire       [15:0]   _zz__19_14_inner_macOut_2;
  reg        [7:0]    _19_14_inner_activation;
  reg        [7:0]    _19_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_14_inner_macOut;

  assign _zz__zz__19_14_inner_macOut = ($signed(io_mulInput) * $signed(_19_14_inner_activation));
  assign _zz__zz__19_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_14_inner_macOut)) ? 16'h007f : _zz__19_14_inner_macOut_2);
  assign _zz__19_14_inner_macOut_2 = (($signed(_zz__19_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_14_inner_activation;
    end else begin
      io_macOut = _19_14_inner_macOut;
    end
  end

  assign _zz__19_14_inner_macOut = ($signed(_zz__zz__19_14_inner_macOut) + $signed(_zz__zz__19_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_14_inner_activation <= 8'h00;
      _19_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_14_inner_activation <= io_addInput;
      end else begin
        _19_14_inner_macOut <= _zz__19_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_621 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_13_inner_macOut;
  wire       [15:0]   _zz__zz__19_13_inner_macOut_1;
  wire       [15:0]   _zz__19_13_inner_macOut_1;
  wire       [15:0]   _zz__19_13_inner_macOut_2;
  reg        [7:0]    _19_13_inner_activation;
  reg        [7:0]    _19_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_13_inner_macOut;

  assign _zz__zz__19_13_inner_macOut = ($signed(io_mulInput) * $signed(_19_13_inner_activation));
  assign _zz__zz__19_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_13_inner_macOut)) ? 16'h007f : _zz__19_13_inner_macOut_2);
  assign _zz__19_13_inner_macOut_2 = (($signed(_zz__19_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_13_inner_activation;
    end else begin
      io_macOut = _19_13_inner_macOut;
    end
  end

  assign _zz__19_13_inner_macOut = ($signed(_zz__zz__19_13_inner_macOut) + $signed(_zz__zz__19_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_13_inner_activation <= 8'h00;
      _19_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_13_inner_activation <= io_addInput;
      end else begin
        _19_13_inner_macOut <= _zz__19_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_620 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_12_inner_macOut;
  wire       [15:0]   _zz__zz__19_12_inner_macOut_1;
  wire       [15:0]   _zz__19_12_inner_macOut_1;
  wire       [15:0]   _zz__19_12_inner_macOut_2;
  reg        [7:0]    _19_12_inner_activation;
  reg        [7:0]    _19_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_12_inner_macOut;

  assign _zz__zz__19_12_inner_macOut = ($signed(io_mulInput) * $signed(_19_12_inner_activation));
  assign _zz__zz__19_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_12_inner_macOut)) ? 16'h007f : _zz__19_12_inner_macOut_2);
  assign _zz__19_12_inner_macOut_2 = (($signed(_zz__19_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_12_inner_activation;
    end else begin
      io_macOut = _19_12_inner_macOut;
    end
  end

  assign _zz__19_12_inner_macOut = ($signed(_zz__zz__19_12_inner_macOut) + $signed(_zz__zz__19_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_12_inner_activation <= 8'h00;
      _19_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_12_inner_activation <= io_addInput;
      end else begin
        _19_12_inner_macOut <= _zz__19_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_619 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_11_inner_macOut;
  wire       [15:0]   _zz__zz__19_11_inner_macOut_1;
  wire       [15:0]   _zz__19_11_inner_macOut_1;
  wire       [15:0]   _zz__19_11_inner_macOut_2;
  reg        [7:0]    _19_11_inner_activation;
  reg        [7:0]    _19_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_11_inner_macOut;

  assign _zz__zz__19_11_inner_macOut = ($signed(io_mulInput) * $signed(_19_11_inner_activation));
  assign _zz__zz__19_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_11_inner_macOut)) ? 16'h007f : _zz__19_11_inner_macOut_2);
  assign _zz__19_11_inner_macOut_2 = (($signed(_zz__19_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_11_inner_activation;
    end else begin
      io_macOut = _19_11_inner_macOut;
    end
  end

  assign _zz__19_11_inner_macOut = ($signed(_zz__zz__19_11_inner_macOut) + $signed(_zz__zz__19_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_11_inner_activation <= 8'h00;
      _19_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_11_inner_activation <= io_addInput;
      end else begin
        _19_11_inner_macOut <= _zz__19_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_618 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_10_inner_macOut;
  wire       [15:0]   _zz__zz__19_10_inner_macOut_1;
  wire       [15:0]   _zz__19_10_inner_macOut_1;
  wire       [15:0]   _zz__19_10_inner_macOut_2;
  reg        [7:0]    _19_10_inner_activation;
  reg        [7:0]    _19_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_10_inner_macOut;

  assign _zz__zz__19_10_inner_macOut = ($signed(io_mulInput) * $signed(_19_10_inner_activation));
  assign _zz__zz__19_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_10_inner_macOut)) ? 16'h007f : _zz__19_10_inner_macOut_2);
  assign _zz__19_10_inner_macOut_2 = (($signed(_zz__19_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_10_inner_activation;
    end else begin
      io_macOut = _19_10_inner_macOut;
    end
  end

  assign _zz__19_10_inner_macOut = ($signed(_zz__zz__19_10_inner_macOut) + $signed(_zz__zz__19_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_10_inner_activation <= 8'h00;
      _19_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_10_inner_activation <= io_addInput;
      end else begin
        _19_10_inner_macOut <= _zz__19_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_617 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_9_inner_macOut;
  wire       [15:0]   _zz__zz__19_9_inner_macOut_1;
  wire       [15:0]   _zz__19_9_inner_macOut_1;
  wire       [15:0]   _zz__19_9_inner_macOut_2;
  reg        [7:0]    _19_9_inner_activation;
  reg        [7:0]    _19_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_9_inner_macOut;

  assign _zz__zz__19_9_inner_macOut = ($signed(io_mulInput) * $signed(_19_9_inner_activation));
  assign _zz__zz__19_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_9_inner_macOut)) ? 16'h007f : _zz__19_9_inner_macOut_2);
  assign _zz__19_9_inner_macOut_2 = (($signed(_zz__19_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_9_inner_activation;
    end else begin
      io_macOut = _19_9_inner_macOut;
    end
  end

  assign _zz__19_9_inner_macOut = ($signed(_zz__zz__19_9_inner_macOut) + $signed(_zz__zz__19_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_9_inner_activation <= 8'h00;
      _19_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_9_inner_activation <= io_addInput;
      end else begin
        _19_9_inner_macOut <= _zz__19_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_616 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_8_inner_macOut;
  wire       [15:0]   _zz__zz__19_8_inner_macOut_1;
  wire       [15:0]   _zz__19_8_inner_macOut_1;
  wire       [15:0]   _zz__19_8_inner_macOut_2;
  reg        [7:0]    _19_8_inner_activation;
  reg        [7:0]    _19_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_8_inner_macOut;

  assign _zz__zz__19_8_inner_macOut = ($signed(io_mulInput) * $signed(_19_8_inner_activation));
  assign _zz__zz__19_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_8_inner_macOut)) ? 16'h007f : _zz__19_8_inner_macOut_2);
  assign _zz__19_8_inner_macOut_2 = (($signed(_zz__19_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_8_inner_activation;
    end else begin
      io_macOut = _19_8_inner_macOut;
    end
  end

  assign _zz__19_8_inner_macOut = ($signed(_zz__zz__19_8_inner_macOut) + $signed(_zz__zz__19_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_8_inner_activation <= 8'h00;
      _19_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_8_inner_activation <= io_addInput;
      end else begin
        _19_8_inner_macOut <= _zz__19_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_615 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_7_inner_macOut;
  wire       [15:0]   _zz__zz__19_7_inner_macOut_1;
  wire       [15:0]   _zz__19_7_inner_macOut_1;
  wire       [15:0]   _zz__19_7_inner_macOut_2;
  reg        [7:0]    _19_7_inner_activation;
  reg        [7:0]    _19_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_7_inner_macOut;

  assign _zz__zz__19_7_inner_macOut = ($signed(io_mulInput) * $signed(_19_7_inner_activation));
  assign _zz__zz__19_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_7_inner_macOut)) ? 16'h007f : _zz__19_7_inner_macOut_2);
  assign _zz__19_7_inner_macOut_2 = (($signed(_zz__19_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_7_inner_activation;
    end else begin
      io_macOut = _19_7_inner_macOut;
    end
  end

  assign _zz__19_7_inner_macOut = ($signed(_zz__zz__19_7_inner_macOut) + $signed(_zz__zz__19_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_7_inner_activation <= 8'h00;
      _19_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_7_inner_activation <= io_addInput;
      end else begin
        _19_7_inner_macOut <= _zz__19_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_614 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_6_inner_macOut;
  wire       [15:0]   _zz__zz__19_6_inner_macOut_1;
  wire       [15:0]   _zz__19_6_inner_macOut_1;
  wire       [15:0]   _zz__19_6_inner_macOut_2;
  reg        [7:0]    _19_6_inner_activation;
  reg        [7:0]    _19_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_6_inner_macOut;

  assign _zz__zz__19_6_inner_macOut = ($signed(io_mulInput) * $signed(_19_6_inner_activation));
  assign _zz__zz__19_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_6_inner_macOut)) ? 16'h007f : _zz__19_6_inner_macOut_2);
  assign _zz__19_6_inner_macOut_2 = (($signed(_zz__19_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_6_inner_activation;
    end else begin
      io_macOut = _19_6_inner_macOut;
    end
  end

  assign _zz__19_6_inner_macOut = ($signed(_zz__zz__19_6_inner_macOut) + $signed(_zz__zz__19_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_6_inner_activation <= 8'h00;
      _19_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_6_inner_activation <= io_addInput;
      end else begin
        _19_6_inner_macOut <= _zz__19_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_613 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_5_inner_macOut;
  wire       [15:0]   _zz__zz__19_5_inner_macOut_1;
  wire       [15:0]   _zz__19_5_inner_macOut_1;
  wire       [15:0]   _zz__19_5_inner_macOut_2;
  reg        [7:0]    _19_5_inner_activation;
  reg        [7:0]    _19_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_5_inner_macOut;

  assign _zz__zz__19_5_inner_macOut = ($signed(io_mulInput) * $signed(_19_5_inner_activation));
  assign _zz__zz__19_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_5_inner_macOut)) ? 16'h007f : _zz__19_5_inner_macOut_2);
  assign _zz__19_5_inner_macOut_2 = (($signed(_zz__19_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_5_inner_activation;
    end else begin
      io_macOut = _19_5_inner_macOut;
    end
  end

  assign _zz__19_5_inner_macOut = ($signed(_zz__zz__19_5_inner_macOut) + $signed(_zz__zz__19_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_5_inner_activation <= 8'h00;
      _19_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_5_inner_activation <= io_addInput;
      end else begin
        _19_5_inner_macOut <= _zz__19_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_612 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_4_inner_macOut;
  wire       [15:0]   _zz__zz__19_4_inner_macOut_1;
  wire       [15:0]   _zz__19_4_inner_macOut_1;
  wire       [15:0]   _zz__19_4_inner_macOut_2;
  reg        [7:0]    _19_4_inner_activation;
  reg        [7:0]    _19_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_4_inner_macOut;

  assign _zz__zz__19_4_inner_macOut = ($signed(io_mulInput) * $signed(_19_4_inner_activation));
  assign _zz__zz__19_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_4_inner_macOut)) ? 16'h007f : _zz__19_4_inner_macOut_2);
  assign _zz__19_4_inner_macOut_2 = (($signed(_zz__19_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_4_inner_activation;
    end else begin
      io_macOut = _19_4_inner_macOut;
    end
  end

  assign _zz__19_4_inner_macOut = ($signed(_zz__zz__19_4_inner_macOut) + $signed(_zz__zz__19_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_4_inner_activation <= 8'h00;
      _19_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_4_inner_activation <= io_addInput;
      end else begin
        _19_4_inner_macOut <= _zz__19_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_611 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_3_inner_macOut;
  wire       [15:0]   _zz__zz__19_3_inner_macOut_1;
  wire       [15:0]   _zz__19_3_inner_macOut_1;
  wire       [15:0]   _zz__19_3_inner_macOut_2;
  reg        [7:0]    _19_3_inner_activation;
  reg        [7:0]    _19_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_3_inner_macOut;

  assign _zz__zz__19_3_inner_macOut = ($signed(io_mulInput) * $signed(_19_3_inner_activation));
  assign _zz__zz__19_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_3_inner_macOut)) ? 16'h007f : _zz__19_3_inner_macOut_2);
  assign _zz__19_3_inner_macOut_2 = (($signed(_zz__19_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_3_inner_activation;
    end else begin
      io_macOut = _19_3_inner_macOut;
    end
  end

  assign _zz__19_3_inner_macOut = ($signed(_zz__zz__19_3_inner_macOut) + $signed(_zz__zz__19_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_3_inner_activation <= 8'h00;
      _19_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_3_inner_activation <= io_addInput;
      end else begin
        _19_3_inner_macOut <= _zz__19_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_610 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_2_inner_macOut;
  wire       [15:0]   _zz__zz__19_2_inner_macOut_1;
  wire       [15:0]   _zz__19_2_inner_macOut_1;
  wire       [15:0]   _zz__19_2_inner_macOut_2;
  reg        [7:0]    _19_2_inner_activation;
  reg        [7:0]    _19_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_2_inner_macOut;

  assign _zz__zz__19_2_inner_macOut = ($signed(io_mulInput) * $signed(_19_2_inner_activation));
  assign _zz__zz__19_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_2_inner_macOut)) ? 16'h007f : _zz__19_2_inner_macOut_2);
  assign _zz__19_2_inner_macOut_2 = (($signed(_zz__19_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_2_inner_activation;
    end else begin
      io_macOut = _19_2_inner_macOut;
    end
  end

  assign _zz__19_2_inner_macOut = ($signed(_zz__zz__19_2_inner_macOut) + $signed(_zz__zz__19_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_2_inner_activation <= 8'h00;
      _19_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_2_inner_activation <= io_addInput;
      end else begin
        _19_2_inner_macOut <= _zz__19_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_609 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_1_inner_macOut;
  wire       [15:0]   _zz__zz__19_1_inner_macOut_1;
  wire       [15:0]   _zz__19_1_inner_macOut_1;
  wire       [15:0]   _zz__19_1_inner_macOut_2;
  reg        [7:0]    _19_1_inner_activation;
  reg        [7:0]    _19_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_1_inner_macOut;

  assign _zz__zz__19_1_inner_macOut = ($signed(io_mulInput) * $signed(_19_1_inner_activation));
  assign _zz__zz__19_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_1_inner_macOut)) ? 16'h007f : _zz__19_1_inner_macOut_2);
  assign _zz__19_1_inner_macOut_2 = (($signed(_zz__19_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_1_inner_activation;
    end else begin
      io_macOut = _19_1_inner_macOut;
    end
  end

  assign _zz__19_1_inner_macOut = ($signed(_zz__zz__19_1_inner_macOut) + $signed(_zz__zz__19_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_1_inner_activation <= 8'h00;
      _19_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_1_inner_activation <= io_addInput;
      end else begin
        _19_1_inner_macOut <= _zz__19_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_608 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__19_0_inner_macOut;
  wire       [15:0]   _zz__zz__19_0_inner_macOut_1;
  wire       [15:0]   _zz__19_0_inner_macOut_1;
  wire       [15:0]   _zz__19_0_inner_macOut_2;
  reg        [7:0]    _19_0_inner_activation;
  reg        [7:0]    _19_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__19_0_inner_macOut;

  assign _zz__zz__19_0_inner_macOut = ($signed(io_mulInput) * $signed(_19_0_inner_activation));
  assign _zz__zz__19_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__19_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__19_0_inner_macOut)) ? 16'h007f : _zz__19_0_inner_macOut_2);
  assign _zz__19_0_inner_macOut_2 = (($signed(_zz__19_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__19_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _19_0_inner_activation;
    end else begin
      io_macOut = _19_0_inner_macOut;
    end
  end

  assign _zz__19_0_inner_macOut = ($signed(_zz__zz__19_0_inner_macOut) + $signed(_zz__zz__19_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _19_0_inner_activation <= 8'h00;
      _19_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _19_0_inner_activation <= io_addInput;
      end else begin
        _19_0_inner_macOut <= _zz__19_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_607 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_31_inner_macOut;
  wire       [15:0]   _zz__zz__18_31_inner_macOut_1;
  wire       [15:0]   _zz__18_31_inner_macOut_1;
  wire       [15:0]   _zz__18_31_inner_macOut_2;
  reg        [7:0]    _18_31_inner_activation;
  reg        [7:0]    _18_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_31_inner_macOut;

  assign _zz__zz__18_31_inner_macOut = ($signed(io_mulInput) * $signed(_18_31_inner_activation));
  assign _zz__zz__18_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_31_inner_macOut)) ? 16'h007f : _zz__18_31_inner_macOut_2);
  assign _zz__18_31_inner_macOut_2 = (($signed(_zz__18_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_31_inner_activation;
    end else begin
      io_macOut = _18_31_inner_macOut;
    end
  end

  assign _zz__18_31_inner_macOut = ($signed(_zz__zz__18_31_inner_macOut) + $signed(_zz__zz__18_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_31_inner_activation <= 8'h00;
      _18_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_31_inner_activation <= io_addInput;
      end else begin
        _18_31_inner_macOut <= _zz__18_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_606 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_30_inner_macOut;
  wire       [15:0]   _zz__zz__18_30_inner_macOut_1;
  wire       [15:0]   _zz__18_30_inner_macOut_1;
  wire       [15:0]   _zz__18_30_inner_macOut_2;
  reg        [7:0]    _18_30_inner_activation;
  reg        [7:0]    _18_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_30_inner_macOut;

  assign _zz__zz__18_30_inner_macOut = ($signed(io_mulInput) * $signed(_18_30_inner_activation));
  assign _zz__zz__18_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_30_inner_macOut)) ? 16'h007f : _zz__18_30_inner_macOut_2);
  assign _zz__18_30_inner_macOut_2 = (($signed(_zz__18_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_30_inner_activation;
    end else begin
      io_macOut = _18_30_inner_macOut;
    end
  end

  assign _zz__18_30_inner_macOut = ($signed(_zz__zz__18_30_inner_macOut) + $signed(_zz__zz__18_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_30_inner_activation <= 8'h00;
      _18_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_30_inner_activation <= io_addInput;
      end else begin
        _18_30_inner_macOut <= _zz__18_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_605 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_29_inner_macOut;
  wire       [15:0]   _zz__zz__18_29_inner_macOut_1;
  wire       [15:0]   _zz__18_29_inner_macOut_1;
  wire       [15:0]   _zz__18_29_inner_macOut_2;
  reg        [7:0]    _18_29_inner_activation;
  reg        [7:0]    _18_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_29_inner_macOut;

  assign _zz__zz__18_29_inner_macOut = ($signed(io_mulInput) * $signed(_18_29_inner_activation));
  assign _zz__zz__18_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_29_inner_macOut)) ? 16'h007f : _zz__18_29_inner_macOut_2);
  assign _zz__18_29_inner_macOut_2 = (($signed(_zz__18_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_29_inner_activation;
    end else begin
      io_macOut = _18_29_inner_macOut;
    end
  end

  assign _zz__18_29_inner_macOut = ($signed(_zz__zz__18_29_inner_macOut) + $signed(_zz__zz__18_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_29_inner_activation <= 8'h00;
      _18_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_29_inner_activation <= io_addInput;
      end else begin
        _18_29_inner_macOut <= _zz__18_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_604 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_28_inner_macOut;
  wire       [15:0]   _zz__zz__18_28_inner_macOut_1;
  wire       [15:0]   _zz__18_28_inner_macOut_1;
  wire       [15:0]   _zz__18_28_inner_macOut_2;
  reg        [7:0]    _18_28_inner_activation;
  reg        [7:0]    _18_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_28_inner_macOut;

  assign _zz__zz__18_28_inner_macOut = ($signed(io_mulInput) * $signed(_18_28_inner_activation));
  assign _zz__zz__18_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_28_inner_macOut)) ? 16'h007f : _zz__18_28_inner_macOut_2);
  assign _zz__18_28_inner_macOut_2 = (($signed(_zz__18_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_28_inner_activation;
    end else begin
      io_macOut = _18_28_inner_macOut;
    end
  end

  assign _zz__18_28_inner_macOut = ($signed(_zz__zz__18_28_inner_macOut) + $signed(_zz__zz__18_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_28_inner_activation <= 8'h00;
      _18_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_28_inner_activation <= io_addInput;
      end else begin
        _18_28_inner_macOut <= _zz__18_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_603 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_27_inner_macOut;
  wire       [15:0]   _zz__zz__18_27_inner_macOut_1;
  wire       [15:0]   _zz__18_27_inner_macOut_1;
  wire       [15:0]   _zz__18_27_inner_macOut_2;
  reg        [7:0]    _18_27_inner_activation;
  reg        [7:0]    _18_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_27_inner_macOut;

  assign _zz__zz__18_27_inner_macOut = ($signed(io_mulInput) * $signed(_18_27_inner_activation));
  assign _zz__zz__18_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_27_inner_macOut)) ? 16'h007f : _zz__18_27_inner_macOut_2);
  assign _zz__18_27_inner_macOut_2 = (($signed(_zz__18_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_27_inner_activation;
    end else begin
      io_macOut = _18_27_inner_macOut;
    end
  end

  assign _zz__18_27_inner_macOut = ($signed(_zz__zz__18_27_inner_macOut) + $signed(_zz__zz__18_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_27_inner_activation <= 8'h00;
      _18_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_27_inner_activation <= io_addInput;
      end else begin
        _18_27_inner_macOut <= _zz__18_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_602 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_26_inner_macOut;
  wire       [15:0]   _zz__zz__18_26_inner_macOut_1;
  wire       [15:0]   _zz__18_26_inner_macOut_1;
  wire       [15:0]   _zz__18_26_inner_macOut_2;
  reg        [7:0]    _18_26_inner_activation;
  reg        [7:0]    _18_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_26_inner_macOut;

  assign _zz__zz__18_26_inner_macOut = ($signed(io_mulInput) * $signed(_18_26_inner_activation));
  assign _zz__zz__18_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_26_inner_macOut)) ? 16'h007f : _zz__18_26_inner_macOut_2);
  assign _zz__18_26_inner_macOut_2 = (($signed(_zz__18_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_26_inner_activation;
    end else begin
      io_macOut = _18_26_inner_macOut;
    end
  end

  assign _zz__18_26_inner_macOut = ($signed(_zz__zz__18_26_inner_macOut) + $signed(_zz__zz__18_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_26_inner_activation <= 8'h00;
      _18_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_26_inner_activation <= io_addInput;
      end else begin
        _18_26_inner_macOut <= _zz__18_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_601 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_25_inner_macOut;
  wire       [15:0]   _zz__zz__18_25_inner_macOut_1;
  wire       [15:0]   _zz__18_25_inner_macOut_1;
  wire       [15:0]   _zz__18_25_inner_macOut_2;
  reg        [7:0]    _18_25_inner_activation;
  reg        [7:0]    _18_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_25_inner_macOut;

  assign _zz__zz__18_25_inner_macOut = ($signed(io_mulInput) * $signed(_18_25_inner_activation));
  assign _zz__zz__18_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_25_inner_macOut)) ? 16'h007f : _zz__18_25_inner_macOut_2);
  assign _zz__18_25_inner_macOut_2 = (($signed(_zz__18_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_25_inner_activation;
    end else begin
      io_macOut = _18_25_inner_macOut;
    end
  end

  assign _zz__18_25_inner_macOut = ($signed(_zz__zz__18_25_inner_macOut) + $signed(_zz__zz__18_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_25_inner_activation <= 8'h00;
      _18_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_25_inner_activation <= io_addInput;
      end else begin
        _18_25_inner_macOut <= _zz__18_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_600 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_24_inner_macOut;
  wire       [15:0]   _zz__zz__18_24_inner_macOut_1;
  wire       [15:0]   _zz__18_24_inner_macOut_1;
  wire       [15:0]   _zz__18_24_inner_macOut_2;
  reg        [7:0]    _18_24_inner_activation;
  reg        [7:0]    _18_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_24_inner_macOut;

  assign _zz__zz__18_24_inner_macOut = ($signed(io_mulInput) * $signed(_18_24_inner_activation));
  assign _zz__zz__18_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_24_inner_macOut)) ? 16'h007f : _zz__18_24_inner_macOut_2);
  assign _zz__18_24_inner_macOut_2 = (($signed(_zz__18_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_24_inner_activation;
    end else begin
      io_macOut = _18_24_inner_macOut;
    end
  end

  assign _zz__18_24_inner_macOut = ($signed(_zz__zz__18_24_inner_macOut) + $signed(_zz__zz__18_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_24_inner_activation <= 8'h00;
      _18_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_24_inner_activation <= io_addInput;
      end else begin
        _18_24_inner_macOut <= _zz__18_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_599 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_23_inner_macOut;
  wire       [15:0]   _zz__zz__18_23_inner_macOut_1;
  wire       [15:0]   _zz__18_23_inner_macOut_1;
  wire       [15:0]   _zz__18_23_inner_macOut_2;
  reg        [7:0]    _18_23_inner_activation;
  reg        [7:0]    _18_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_23_inner_macOut;

  assign _zz__zz__18_23_inner_macOut = ($signed(io_mulInput) * $signed(_18_23_inner_activation));
  assign _zz__zz__18_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_23_inner_macOut)) ? 16'h007f : _zz__18_23_inner_macOut_2);
  assign _zz__18_23_inner_macOut_2 = (($signed(_zz__18_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_23_inner_activation;
    end else begin
      io_macOut = _18_23_inner_macOut;
    end
  end

  assign _zz__18_23_inner_macOut = ($signed(_zz__zz__18_23_inner_macOut) + $signed(_zz__zz__18_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_23_inner_activation <= 8'h00;
      _18_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_23_inner_activation <= io_addInput;
      end else begin
        _18_23_inner_macOut <= _zz__18_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_598 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_22_inner_macOut;
  wire       [15:0]   _zz__zz__18_22_inner_macOut_1;
  wire       [15:0]   _zz__18_22_inner_macOut_1;
  wire       [15:0]   _zz__18_22_inner_macOut_2;
  reg        [7:0]    _18_22_inner_activation;
  reg        [7:0]    _18_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_22_inner_macOut;

  assign _zz__zz__18_22_inner_macOut = ($signed(io_mulInput) * $signed(_18_22_inner_activation));
  assign _zz__zz__18_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_22_inner_macOut)) ? 16'h007f : _zz__18_22_inner_macOut_2);
  assign _zz__18_22_inner_macOut_2 = (($signed(_zz__18_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_22_inner_activation;
    end else begin
      io_macOut = _18_22_inner_macOut;
    end
  end

  assign _zz__18_22_inner_macOut = ($signed(_zz__zz__18_22_inner_macOut) + $signed(_zz__zz__18_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_22_inner_activation <= 8'h00;
      _18_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_22_inner_activation <= io_addInput;
      end else begin
        _18_22_inner_macOut <= _zz__18_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_597 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_21_inner_macOut;
  wire       [15:0]   _zz__zz__18_21_inner_macOut_1;
  wire       [15:0]   _zz__18_21_inner_macOut_1;
  wire       [15:0]   _zz__18_21_inner_macOut_2;
  reg        [7:0]    _18_21_inner_activation;
  reg        [7:0]    _18_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_21_inner_macOut;

  assign _zz__zz__18_21_inner_macOut = ($signed(io_mulInput) * $signed(_18_21_inner_activation));
  assign _zz__zz__18_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_21_inner_macOut)) ? 16'h007f : _zz__18_21_inner_macOut_2);
  assign _zz__18_21_inner_macOut_2 = (($signed(_zz__18_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_21_inner_activation;
    end else begin
      io_macOut = _18_21_inner_macOut;
    end
  end

  assign _zz__18_21_inner_macOut = ($signed(_zz__zz__18_21_inner_macOut) + $signed(_zz__zz__18_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_21_inner_activation <= 8'h00;
      _18_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_21_inner_activation <= io_addInput;
      end else begin
        _18_21_inner_macOut <= _zz__18_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_596 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_20_inner_macOut;
  wire       [15:0]   _zz__zz__18_20_inner_macOut_1;
  wire       [15:0]   _zz__18_20_inner_macOut_1;
  wire       [15:0]   _zz__18_20_inner_macOut_2;
  reg        [7:0]    _18_20_inner_activation;
  reg        [7:0]    _18_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_20_inner_macOut;

  assign _zz__zz__18_20_inner_macOut = ($signed(io_mulInput) * $signed(_18_20_inner_activation));
  assign _zz__zz__18_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_20_inner_macOut)) ? 16'h007f : _zz__18_20_inner_macOut_2);
  assign _zz__18_20_inner_macOut_2 = (($signed(_zz__18_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_20_inner_activation;
    end else begin
      io_macOut = _18_20_inner_macOut;
    end
  end

  assign _zz__18_20_inner_macOut = ($signed(_zz__zz__18_20_inner_macOut) + $signed(_zz__zz__18_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_20_inner_activation <= 8'h00;
      _18_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_20_inner_activation <= io_addInput;
      end else begin
        _18_20_inner_macOut <= _zz__18_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_595 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_19_inner_macOut;
  wire       [15:0]   _zz__zz__18_19_inner_macOut_1;
  wire       [15:0]   _zz__18_19_inner_macOut_1;
  wire       [15:0]   _zz__18_19_inner_macOut_2;
  reg        [7:0]    _18_19_inner_activation;
  reg        [7:0]    _18_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_19_inner_macOut;

  assign _zz__zz__18_19_inner_macOut = ($signed(io_mulInput) * $signed(_18_19_inner_activation));
  assign _zz__zz__18_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_19_inner_macOut)) ? 16'h007f : _zz__18_19_inner_macOut_2);
  assign _zz__18_19_inner_macOut_2 = (($signed(_zz__18_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_19_inner_activation;
    end else begin
      io_macOut = _18_19_inner_macOut;
    end
  end

  assign _zz__18_19_inner_macOut = ($signed(_zz__zz__18_19_inner_macOut) + $signed(_zz__zz__18_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_19_inner_activation <= 8'h00;
      _18_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_19_inner_activation <= io_addInput;
      end else begin
        _18_19_inner_macOut <= _zz__18_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_594 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_18_inner_macOut;
  wire       [15:0]   _zz__zz__18_18_inner_macOut_1;
  wire       [15:0]   _zz__18_18_inner_macOut_1;
  wire       [15:0]   _zz__18_18_inner_macOut_2;
  reg        [7:0]    _18_18_inner_activation;
  reg        [7:0]    _18_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_18_inner_macOut;

  assign _zz__zz__18_18_inner_macOut = ($signed(io_mulInput) * $signed(_18_18_inner_activation));
  assign _zz__zz__18_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_18_inner_macOut)) ? 16'h007f : _zz__18_18_inner_macOut_2);
  assign _zz__18_18_inner_macOut_2 = (($signed(_zz__18_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_18_inner_activation;
    end else begin
      io_macOut = _18_18_inner_macOut;
    end
  end

  assign _zz__18_18_inner_macOut = ($signed(_zz__zz__18_18_inner_macOut) + $signed(_zz__zz__18_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_18_inner_activation <= 8'h00;
      _18_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_18_inner_activation <= io_addInput;
      end else begin
        _18_18_inner_macOut <= _zz__18_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_593 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_17_inner_macOut;
  wire       [15:0]   _zz__zz__18_17_inner_macOut_1;
  wire       [15:0]   _zz__18_17_inner_macOut_1;
  wire       [15:0]   _zz__18_17_inner_macOut_2;
  reg        [7:0]    _18_17_inner_activation;
  reg        [7:0]    _18_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_17_inner_macOut;

  assign _zz__zz__18_17_inner_macOut = ($signed(io_mulInput) * $signed(_18_17_inner_activation));
  assign _zz__zz__18_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_17_inner_macOut)) ? 16'h007f : _zz__18_17_inner_macOut_2);
  assign _zz__18_17_inner_macOut_2 = (($signed(_zz__18_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_17_inner_activation;
    end else begin
      io_macOut = _18_17_inner_macOut;
    end
  end

  assign _zz__18_17_inner_macOut = ($signed(_zz__zz__18_17_inner_macOut) + $signed(_zz__zz__18_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_17_inner_activation <= 8'h00;
      _18_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_17_inner_activation <= io_addInput;
      end else begin
        _18_17_inner_macOut <= _zz__18_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_592 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_16_inner_macOut;
  wire       [15:0]   _zz__zz__18_16_inner_macOut_1;
  wire       [15:0]   _zz__18_16_inner_macOut_1;
  wire       [15:0]   _zz__18_16_inner_macOut_2;
  reg        [7:0]    _18_16_inner_activation;
  reg        [7:0]    _18_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_16_inner_macOut;

  assign _zz__zz__18_16_inner_macOut = ($signed(io_mulInput) * $signed(_18_16_inner_activation));
  assign _zz__zz__18_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_16_inner_macOut)) ? 16'h007f : _zz__18_16_inner_macOut_2);
  assign _zz__18_16_inner_macOut_2 = (($signed(_zz__18_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_16_inner_activation;
    end else begin
      io_macOut = _18_16_inner_macOut;
    end
  end

  assign _zz__18_16_inner_macOut = ($signed(_zz__zz__18_16_inner_macOut) + $signed(_zz__zz__18_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_16_inner_activation <= 8'h00;
      _18_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_16_inner_activation <= io_addInput;
      end else begin
        _18_16_inner_macOut <= _zz__18_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_591 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_15_inner_macOut;
  wire       [15:0]   _zz__zz__18_15_inner_macOut_1;
  wire       [15:0]   _zz__18_15_inner_macOut_1;
  wire       [15:0]   _zz__18_15_inner_macOut_2;
  reg        [7:0]    _18_15_inner_activation;
  reg        [7:0]    _18_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_15_inner_macOut;

  assign _zz__zz__18_15_inner_macOut = ($signed(io_mulInput) * $signed(_18_15_inner_activation));
  assign _zz__zz__18_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_15_inner_macOut)) ? 16'h007f : _zz__18_15_inner_macOut_2);
  assign _zz__18_15_inner_macOut_2 = (($signed(_zz__18_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_15_inner_activation;
    end else begin
      io_macOut = _18_15_inner_macOut;
    end
  end

  assign _zz__18_15_inner_macOut = ($signed(_zz__zz__18_15_inner_macOut) + $signed(_zz__zz__18_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_15_inner_activation <= 8'h00;
      _18_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_15_inner_activation <= io_addInput;
      end else begin
        _18_15_inner_macOut <= _zz__18_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_590 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_14_inner_macOut;
  wire       [15:0]   _zz__zz__18_14_inner_macOut_1;
  wire       [15:0]   _zz__18_14_inner_macOut_1;
  wire       [15:0]   _zz__18_14_inner_macOut_2;
  reg        [7:0]    _18_14_inner_activation;
  reg        [7:0]    _18_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_14_inner_macOut;

  assign _zz__zz__18_14_inner_macOut = ($signed(io_mulInput) * $signed(_18_14_inner_activation));
  assign _zz__zz__18_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_14_inner_macOut)) ? 16'h007f : _zz__18_14_inner_macOut_2);
  assign _zz__18_14_inner_macOut_2 = (($signed(_zz__18_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_14_inner_activation;
    end else begin
      io_macOut = _18_14_inner_macOut;
    end
  end

  assign _zz__18_14_inner_macOut = ($signed(_zz__zz__18_14_inner_macOut) + $signed(_zz__zz__18_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_14_inner_activation <= 8'h00;
      _18_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_14_inner_activation <= io_addInput;
      end else begin
        _18_14_inner_macOut <= _zz__18_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_589 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_13_inner_macOut;
  wire       [15:0]   _zz__zz__18_13_inner_macOut_1;
  wire       [15:0]   _zz__18_13_inner_macOut_1;
  wire       [15:0]   _zz__18_13_inner_macOut_2;
  reg        [7:0]    _18_13_inner_activation;
  reg        [7:0]    _18_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_13_inner_macOut;

  assign _zz__zz__18_13_inner_macOut = ($signed(io_mulInput) * $signed(_18_13_inner_activation));
  assign _zz__zz__18_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_13_inner_macOut)) ? 16'h007f : _zz__18_13_inner_macOut_2);
  assign _zz__18_13_inner_macOut_2 = (($signed(_zz__18_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_13_inner_activation;
    end else begin
      io_macOut = _18_13_inner_macOut;
    end
  end

  assign _zz__18_13_inner_macOut = ($signed(_zz__zz__18_13_inner_macOut) + $signed(_zz__zz__18_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_13_inner_activation <= 8'h00;
      _18_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_13_inner_activation <= io_addInput;
      end else begin
        _18_13_inner_macOut <= _zz__18_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_588 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_12_inner_macOut;
  wire       [15:0]   _zz__zz__18_12_inner_macOut_1;
  wire       [15:0]   _zz__18_12_inner_macOut_1;
  wire       [15:0]   _zz__18_12_inner_macOut_2;
  reg        [7:0]    _18_12_inner_activation;
  reg        [7:0]    _18_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_12_inner_macOut;

  assign _zz__zz__18_12_inner_macOut = ($signed(io_mulInput) * $signed(_18_12_inner_activation));
  assign _zz__zz__18_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_12_inner_macOut)) ? 16'h007f : _zz__18_12_inner_macOut_2);
  assign _zz__18_12_inner_macOut_2 = (($signed(_zz__18_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_12_inner_activation;
    end else begin
      io_macOut = _18_12_inner_macOut;
    end
  end

  assign _zz__18_12_inner_macOut = ($signed(_zz__zz__18_12_inner_macOut) + $signed(_zz__zz__18_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_12_inner_activation <= 8'h00;
      _18_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_12_inner_activation <= io_addInput;
      end else begin
        _18_12_inner_macOut <= _zz__18_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_587 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_11_inner_macOut;
  wire       [15:0]   _zz__zz__18_11_inner_macOut_1;
  wire       [15:0]   _zz__18_11_inner_macOut_1;
  wire       [15:0]   _zz__18_11_inner_macOut_2;
  reg        [7:0]    _18_11_inner_activation;
  reg        [7:0]    _18_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_11_inner_macOut;

  assign _zz__zz__18_11_inner_macOut = ($signed(io_mulInput) * $signed(_18_11_inner_activation));
  assign _zz__zz__18_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_11_inner_macOut)) ? 16'h007f : _zz__18_11_inner_macOut_2);
  assign _zz__18_11_inner_macOut_2 = (($signed(_zz__18_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_11_inner_activation;
    end else begin
      io_macOut = _18_11_inner_macOut;
    end
  end

  assign _zz__18_11_inner_macOut = ($signed(_zz__zz__18_11_inner_macOut) + $signed(_zz__zz__18_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_11_inner_activation <= 8'h00;
      _18_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_11_inner_activation <= io_addInput;
      end else begin
        _18_11_inner_macOut <= _zz__18_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_586 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_10_inner_macOut;
  wire       [15:0]   _zz__zz__18_10_inner_macOut_1;
  wire       [15:0]   _zz__18_10_inner_macOut_1;
  wire       [15:0]   _zz__18_10_inner_macOut_2;
  reg        [7:0]    _18_10_inner_activation;
  reg        [7:0]    _18_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_10_inner_macOut;

  assign _zz__zz__18_10_inner_macOut = ($signed(io_mulInput) * $signed(_18_10_inner_activation));
  assign _zz__zz__18_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_10_inner_macOut)) ? 16'h007f : _zz__18_10_inner_macOut_2);
  assign _zz__18_10_inner_macOut_2 = (($signed(_zz__18_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_10_inner_activation;
    end else begin
      io_macOut = _18_10_inner_macOut;
    end
  end

  assign _zz__18_10_inner_macOut = ($signed(_zz__zz__18_10_inner_macOut) + $signed(_zz__zz__18_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_10_inner_activation <= 8'h00;
      _18_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_10_inner_activation <= io_addInput;
      end else begin
        _18_10_inner_macOut <= _zz__18_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_585 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_9_inner_macOut;
  wire       [15:0]   _zz__zz__18_9_inner_macOut_1;
  wire       [15:0]   _zz__18_9_inner_macOut_1;
  wire       [15:0]   _zz__18_9_inner_macOut_2;
  reg        [7:0]    _18_9_inner_activation;
  reg        [7:0]    _18_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_9_inner_macOut;

  assign _zz__zz__18_9_inner_macOut = ($signed(io_mulInput) * $signed(_18_9_inner_activation));
  assign _zz__zz__18_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_9_inner_macOut)) ? 16'h007f : _zz__18_9_inner_macOut_2);
  assign _zz__18_9_inner_macOut_2 = (($signed(_zz__18_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_9_inner_activation;
    end else begin
      io_macOut = _18_9_inner_macOut;
    end
  end

  assign _zz__18_9_inner_macOut = ($signed(_zz__zz__18_9_inner_macOut) + $signed(_zz__zz__18_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_9_inner_activation <= 8'h00;
      _18_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_9_inner_activation <= io_addInput;
      end else begin
        _18_9_inner_macOut <= _zz__18_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_584 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_8_inner_macOut;
  wire       [15:0]   _zz__zz__18_8_inner_macOut_1;
  wire       [15:0]   _zz__18_8_inner_macOut_1;
  wire       [15:0]   _zz__18_8_inner_macOut_2;
  reg        [7:0]    _18_8_inner_activation;
  reg        [7:0]    _18_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_8_inner_macOut;

  assign _zz__zz__18_8_inner_macOut = ($signed(io_mulInput) * $signed(_18_8_inner_activation));
  assign _zz__zz__18_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_8_inner_macOut)) ? 16'h007f : _zz__18_8_inner_macOut_2);
  assign _zz__18_8_inner_macOut_2 = (($signed(_zz__18_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_8_inner_activation;
    end else begin
      io_macOut = _18_8_inner_macOut;
    end
  end

  assign _zz__18_8_inner_macOut = ($signed(_zz__zz__18_8_inner_macOut) + $signed(_zz__zz__18_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_8_inner_activation <= 8'h00;
      _18_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_8_inner_activation <= io_addInput;
      end else begin
        _18_8_inner_macOut <= _zz__18_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_583 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_7_inner_macOut;
  wire       [15:0]   _zz__zz__18_7_inner_macOut_1;
  wire       [15:0]   _zz__18_7_inner_macOut_1;
  wire       [15:0]   _zz__18_7_inner_macOut_2;
  reg        [7:0]    _18_7_inner_activation;
  reg        [7:0]    _18_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_7_inner_macOut;

  assign _zz__zz__18_7_inner_macOut = ($signed(io_mulInput) * $signed(_18_7_inner_activation));
  assign _zz__zz__18_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_7_inner_macOut)) ? 16'h007f : _zz__18_7_inner_macOut_2);
  assign _zz__18_7_inner_macOut_2 = (($signed(_zz__18_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_7_inner_activation;
    end else begin
      io_macOut = _18_7_inner_macOut;
    end
  end

  assign _zz__18_7_inner_macOut = ($signed(_zz__zz__18_7_inner_macOut) + $signed(_zz__zz__18_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_7_inner_activation <= 8'h00;
      _18_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_7_inner_activation <= io_addInput;
      end else begin
        _18_7_inner_macOut <= _zz__18_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_582 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_6_inner_macOut;
  wire       [15:0]   _zz__zz__18_6_inner_macOut_1;
  wire       [15:0]   _zz__18_6_inner_macOut_1;
  wire       [15:0]   _zz__18_6_inner_macOut_2;
  reg        [7:0]    _18_6_inner_activation;
  reg        [7:0]    _18_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_6_inner_macOut;

  assign _zz__zz__18_6_inner_macOut = ($signed(io_mulInput) * $signed(_18_6_inner_activation));
  assign _zz__zz__18_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_6_inner_macOut)) ? 16'h007f : _zz__18_6_inner_macOut_2);
  assign _zz__18_6_inner_macOut_2 = (($signed(_zz__18_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_6_inner_activation;
    end else begin
      io_macOut = _18_6_inner_macOut;
    end
  end

  assign _zz__18_6_inner_macOut = ($signed(_zz__zz__18_6_inner_macOut) + $signed(_zz__zz__18_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_6_inner_activation <= 8'h00;
      _18_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_6_inner_activation <= io_addInput;
      end else begin
        _18_6_inner_macOut <= _zz__18_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_581 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_5_inner_macOut;
  wire       [15:0]   _zz__zz__18_5_inner_macOut_1;
  wire       [15:0]   _zz__18_5_inner_macOut_1;
  wire       [15:0]   _zz__18_5_inner_macOut_2;
  reg        [7:0]    _18_5_inner_activation;
  reg        [7:0]    _18_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_5_inner_macOut;

  assign _zz__zz__18_5_inner_macOut = ($signed(io_mulInput) * $signed(_18_5_inner_activation));
  assign _zz__zz__18_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_5_inner_macOut)) ? 16'h007f : _zz__18_5_inner_macOut_2);
  assign _zz__18_5_inner_macOut_2 = (($signed(_zz__18_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_5_inner_activation;
    end else begin
      io_macOut = _18_5_inner_macOut;
    end
  end

  assign _zz__18_5_inner_macOut = ($signed(_zz__zz__18_5_inner_macOut) + $signed(_zz__zz__18_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_5_inner_activation <= 8'h00;
      _18_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_5_inner_activation <= io_addInput;
      end else begin
        _18_5_inner_macOut <= _zz__18_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_580 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_4_inner_macOut;
  wire       [15:0]   _zz__zz__18_4_inner_macOut_1;
  wire       [15:0]   _zz__18_4_inner_macOut_1;
  wire       [15:0]   _zz__18_4_inner_macOut_2;
  reg        [7:0]    _18_4_inner_activation;
  reg        [7:0]    _18_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_4_inner_macOut;

  assign _zz__zz__18_4_inner_macOut = ($signed(io_mulInput) * $signed(_18_4_inner_activation));
  assign _zz__zz__18_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_4_inner_macOut)) ? 16'h007f : _zz__18_4_inner_macOut_2);
  assign _zz__18_4_inner_macOut_2 = (($signed(_zz__18_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_4_inner_activation;
    end else begin
      io_macOut = _18_4_inner_macOut;
    end
  end

  assign _zz__18_4_inner_macOut = ($signed(_zz__zz__18_4_inner_macOut) + $signed(_zz__zz__18_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_4_inner_activation <= 8'h00;
      _18_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_4_inner_activation <= io_addInput;
      end else begin
        _18_4_inner_macOut <= _zz__18_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_579 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_3_inner_macOut;
  wire       [15:0]   _zz__zz__18_3_inner_macOut_1;
  wire       [15:0]   _zz__18_3_inner_macOut_1;
  wire       [15:0]   _zz__18_3_inner_macOut_2;
  reg        [7:0]    _18_3_inner_activation;
  reg        [7:0]    _18_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_3_inner_macOut;

  assign _zz__zz__18_3_inner_macOut = ($signed(io_mulInput) * $signed(_18_3_inner_activation));
  assign _zz__zz__18_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_3_inner_macOut)) ? 16'h007f : _zz__18_3_inner_macOut_2);
  assign _zz__18_3_inner_macOut_2 = (($signed(_zz__18_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_3_inner_activation;
    end else begin
      io_macOut = _18_3_inner_macOut;
    end
  end

  assign _zz__18_3_inner_macOut = ($signed(_zz__zz__18_3_inner_macOut) + $signed(_zz__zz__18_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_3_inner_activation <= 8'h00;
      _18_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_3_inner_activation <= io_addInput;
      end else begin
        _18_3_inner_macOut <= _zz__18_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_578 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_2_inner_macOut;
  wire       [15:0]   _zz__zz__18_2_inner_macOut_1;
  wire       [15:0]   _zz__18_2_inner_macOut_1;
  wire       [15:0]   _zz__18_2_inner_macOut_2;
  reg        [7:0]    _18_2_inner_activation;
  reg        [7:0]    _18_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_2_inner_macOut;

  assign _zz__zz__18_2_inner_macOut = ($signed(io_mulInput) * $signed(_18_2_inner_activation));
  assign _zz__zz__18_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_2_inner_macOut)) ? 16'h007f : _zz__18_2_inner_macOut_2);
  assign _zz__18_2_inner_macOut_2 = (($signed(_zz__18_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_2_inner_activation;
    end else begin
      io_macOut = _18_2_inner_macOut;
    end
  end

  assign _zz__18_2_inner_macOut = ($signed(_zz__zz__18_2_inner_macOut) + $signed(_zz__zz__18_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_2_inner_activation <= 8'h00;
      _18_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_2_inner_activation <= io_addInput;
      end else begin
        _18_2_inner_macOut <= _zz__18_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_577 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_1_inner_macOut;
  wire       [15:0]   _zz__zz__18_1_inner_macOut_1;
  wire       [15:0]   _zz__18_1_inner_macOut_1;
  wire       [15:0]   _zz__18_1_inner_macOut_2;
  reg        [7:0]    _18_1_inner_activation;
  reg        [7:0]    _18_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_1_inner_macOut;

  assign _zz__zz__18_1_inner_macOut = ($signed(io_mulInput) * $signed(_18_1_inner_activation));
  assign _zz__zz__18_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_1_inner_macOut)) ? 16'h007f : _zz__18_1_inner_macOut_2);
  assign _zz__18_1_inner_macOut_2 = (($signed(_zz__18_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_1_inner_activation;
    end else begin
      io_macOut = _18_1_inner_macOut;
    end
  end

  assign _zz__18_1_inner_macOut = ($signed(_zz__zz__18_1_inner_macOut) + $signed(_zz__zz__18_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_1_inner_activation <= 8'h00;
      _18_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_1_inner_activation <= io_addInput;
      end else begin
        _18_1_inner_macOut <= _zz__18_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_576 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__18_0_inner_macOut;
  wire       [15:0]   _zz__zz__18_0_inner_macOut_1;
  wire       [15:0]   _zz__18_0_inner_macOut_1;
  wire       [15:0]   _zz__18_0_inner_macOut_2;
  reg        [7:0]    _18_0_inner_activation;
  reg        [7:0]    _18_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__18_0_inner_macOut;

  assign _zz__zz__18_0_inner_macOut = ($signed(io_mulInput) * $signed(_18_0_inner_activation));
  assign _zz__zz__18_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__18_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__18_0_inner_macOut)) ? 16'h007f : _zz__18_0_inner_macOut_2);
  assign _zz__18_0_inner_macOut_2 = (($signed(_zz__18_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__18_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _18_0_inner_activation;
    end else begin
      io_macOut = _18_0_inner_macOut;
    end
  end

  assign _zz__18_0_inner_macOut = ($signed(_zz__zz__18_0_inner_macOut) + $signed(_zz__zz__18_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _18_0_inner_activation <= 8'h00;
      _18_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _18_0_inner_activation <= io_addInput;
      end else begin
        _18_0_inner_macOut <= _zz__18_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_575 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_31_inner_macOut;
  wire       [15:0]   _zz__zz__17_31_inner_macOut_1;
  wire       [15:0]   _zz__17_31_inner_macOut_1;
  wire       [15:0]   _zz__17_31_inner_macOut_2;
  reg        [7:0]    _17_31_inner_activation;
  reg        [7:0]    _17_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_31_inner_macOut;

  assign _zz__zz__17_31_inner_macOut = ($signed(io_mulInput) * $signed(_17_31_inner_activation));
  assign _zz__zz__17_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_31_inner_macOut)) ? 16'h007f : _zz__17_31_inner_macOut_2);
  assign _zz__17_31_inner_macOut_2 = (($signed(_zz__17_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_31_inner_activation;
    end else begin
      io_macOut = _17_31_inner_macOut;
    end
  end

  assign _zz__17_31_inner_macOut = ($signed(_zz__zz__17_31_inner_macOut) + $signed(_zz__zz__17_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_31_inner_activation <= 8'h00;
      _17_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_31_inner_activation <= io_addInput;
      end else begin
        _17_31_inner_macOut <= _zz__17_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_574 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_30_inner_macOut;
  wire       [15:0]   _zz__zz__17_30_inner_macOut_1;
  wire       [15:0]   _zz__17_30_inner_macOut_1;
  wire       [15:0]   _zz__17_30_inner_macOut_2;
  reg        [7:0]    _17_30_inner_activation;
  reg        [7:0]    _17_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_30_inner_macOut;

  assign _zz__zz__17_30_inner_macOut = ($signed(io_mulInput) * $signed(_17_30_inner_activation));
  assign _zz__zz__17_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_30_inner_macOut)) ? 16'h007f : _zz__17_30_inner_macOut_2);
  assign _zz__17_30_inner_macOut_2 = (($signed(_zz__17_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_30_inner_activation;
    end else begin
      io_macOut = _17_30_inner_macOut;
    end
  end

  assign _zz__17_30_inner_macOut = ($signed(_zz__zz__17_30_inner_macOut) + $signed(_zz__zz__17_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_30_inner_activation <= 8'h00;
      _17_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_30_inner_activation <= io_addInput;
      end else begin
        _17_30_inner_macOut <= _zz__17_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_573 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_29_inner_macOut;
  wire       [15:0]   _zz__zz__17_29_inner_macOut_1;
  wire       [15:0]   _zz__17_29_inner_macOut_1;
  wire       [15:0]   _zz__17_29_inner_macOut_2;
  reg        [7:0]    _17_29_inner_activation;
  reg        [7:0]    _17_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_29_inner_macOut;

  assign _zz__zz__17_29_inner_macOut = ($signed(io_mulInput) * $signed(_17_29_inner_activation));
  assign _zz__zz__17_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_29_inner_macOut)) ? 16'h007f : _zz__17_29_inner_macOut_2);
  assign _zz__17_29_inner_macOut_2 = (($signed(_zz__17_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_29_inner_activation;
    end else begin
      io_macOut = _17_29_inner_macOut;
    end
  end

  assign _zz__17_29_inner_macOut = ($signed(_zz__zz__17_29_inner_macOut) + $signed(_zz__zz__17_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_29_inner_activation <= 8'h00;
      _17_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_29_inner_activation <= io_addInput;
      end else begin
        _17_29_inner_macOut <= _zz__17_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_572 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_28_inner_macOut;
  wire       [15:0]   _zz__zz__17_28_inner_macOut_1;
  wire       [15:0]   _zz__17_28_inner_macOut_1;
  wire       [15:0]   _zz__17_28_inner_macOut_2;
  reg        [7:0]    _17_28_inner_activation;
  reg        [7:0]    _17_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_28_inner_macOut;

  assign _zz__zz__17_28_inner_macOut = ($signed(io_mulInput) * $signed(_17_28_inner_activation));
  assign _zz__zz__17_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_28_inner_macOut)) ? 16'h007f : _zz__17_28_inner_macOut_2);
  assign _zz__17_28_inner_macOut_2 = (($signed(_zz__17_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_28_inner_activation;
    end else begin
      io_macOut = _17_28_inner_macOut;
    end
  end

  assign _zz__17_28_inner_macOut = ($signed(_zz__zz__17_28_inner_macOut) + $signed(_zz__zz__17_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_28_inner_activation <= 8'h00;
      _17_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_28_inner_activation <= io_addInput;
      end else begin
        _17_28_inner_macOut <= _zz__17_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_571 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_27_inner_macOut;
  wire       [15:0]   _zz__zz__17_27_inner_macOut_1;
  wire       [15:0]   _zz__17_27_inner_macOut_1;
  wire       [15:0]   _zz__17_27_inner_macOut_2;
  reg        [7:0]    _17_27_inner_activation;
  reg        [7:0]    _17_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_27_inner_macOut;

  assign _zz__zz__17_27_inner_macOut = ($signed(io_mulInput) * $signed(_17_27_inner_activation));
  assign _zz__zz__17_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_27_inner_macOut)) ? 16'h007f : _zz__17_27_inner_macOut_2);
  assign _zz__17_27_inner_macOut_2 = (($signed(_zz__17_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_27_inner_activation;
    end else begin
      io_macOut = _17_27_inner_macOut;
    end
  end

  assign _zz__17_27_inner_macOut = ($signed(_zz__zz__17_27_inner_macOut) + $signed(_zz__zz__17_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_27_inner_activation <= 8'h00;
      _17_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_27_inner_activation <= io_addInput;
      end else begin
        _17_27_inner_macOut <= _zz__17_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_570 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_26_inner_macOut;
  wire       [15:0]   _zz__zz__17_26_inner_macOut_1;
  wire       [15:0]   _zz__17_26_inner_macOut_1;
  wire       [15:0]   _zz__17_26_inner_macOut_2;
  reg        [7:0]    _17_26_inner_activation;
  reg        [7:0]    _17_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_26_inner_macOut;

  assign _zz__zz__17_26_inner_macOut = ($signed(io_mulInput) * $signed(_17_26_inner_activation));
  assign _zz__zz__17_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_26_inner_macOut)) ? 16'h007f : _zz__17_26_inner_macOut_2);
  assign _zz__17_26_inner_macOut_2 = (($signed(_zz__17_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_26_inner_activation;
    end else begin
      io_macOut = _17_26_inner_macOut;
    end
  end

  assign _zz__17_26_inner_macOut = ($signed(_zz__zz__17_26_inner_macOut) + $signed(_zz__zz__17_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_26_inner_activation <= 8'h00;
      _17_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_26_inner_activation <= io_addInput;
      end else begin
        _17_26_inner_macOut <= _zz__17_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_569 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_25_inner_macOut;
  wire       [15:0]   _zz__zz__17_25_inner_macOut_1;
  wire       [15:0]   _zz__17_25_inner_macOut_1;
  wire       [15:0]   _zz__17_25_inner_macOut_2;
  reg        [7:0]    _17_25_inner_activation;
  reg        [7:0]    _17_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_25_inner_macOut;

  assign _zz__zz__17_25_inner_macOut = ($signed(io_mulInput) * $signed(_17_25_inner_activation));
  assign _zz__zz__17_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_25_inner_macOut)) ? 16'h007f : _zz__17_25_inner_macOut_2);
  assign _zz__17_25_inner_macOut_2 = (($signed(_zz__17_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_25_inner_activation;
    end else begin
      io_macOut = _17_25_inner_macOut;
    end
  end

  assign _zz__17_25_inner_macOut = ($signed(_zz__zz__17_25_inner_macOut) + $signed(_zz__zz__17_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_25_inner_activation <= 8'h00;
      _17_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_25_inner_activation <= io_addInput;
      end else begin
        _17_25_inner_macOut <= _zz__17_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_568 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_24_inner_macOut;
  wire       [15:0]   _zz__zz__17_24_inner_macOut_1;
  wire       [15:0]   _zz__17_24_inner_macOut_1;
  wire       [15:0]   _zz__17_24_inner_macOut_2;
  reg        [7:0]    _17_24_inner_activation;
  reg        [7:0]    _17_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_24_inner_macOut;

  assign _zz__zz__17_24_inner_macOut = ($signed(io_mulInput) * $signed(_17_24_inner_activation));
  assign _zz__zz__17_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_24_inner_macOut)) ? 16'h007f : _zz__17_24_inner_macOut_2);
  assign _zz__17_24_inner_macOut_2 = (($signed(_zz__17_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_24_inner_activation;
    end else begin
      io_macOut = _17_24_inner_macOut;
    end
  end

  assign _zz__17_24_inner_macOut = ($signed(_zz__zz__17_24_inner_macOut) + $signed(_zz__zz__17_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_24_inner_activation <= 8'h00;
      _17_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_24_inner_activation <= io_addInput;
      end else begin
        _17_24_inner_macOut <= _zz__17_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_567 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_23_inner_macOut;
  wire       [15:0]   _zz__zz__17_23_inner_macOut_1;
  wire       [15:0]   _zz__17_23_inner_macOut_1;
  wire       [15:0]   _zz__17_23_inner_macOut_2;
  reg        [7:0]    _17_23_inner_activation;
  reg        [7:0]    _17_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_23_inner_macOut;

  assign _zz__zz__17_23_inner_macOut = ($signed(io_mulInput) * $signed(_17_23_inner_activation));
  assign _zz__zz__17_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_23_inner_macOut)) ? 16'h007f : _zz__17_23_inner_macOut_2);
  assign _zz__17_23_inner_macOut_2 = (($signed(_zz__17_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_23_inner_activation;
    end else begin
      io_macOut = _17_23_inner_macOut;
    end
  end

  assign _zz__17_23_inner_macOut = ($signed(_zz__zz__17_23_inner_macOut) + $signed(_zz__zz__17_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_23_inner_activation <= 8'h00;
      _17_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_23_inner_activation <= io_addInput;
      end else begin
        _17_23_inner_macOut <= _zz__17_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_566 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_22_inner_macOut;
  wire       [15:0]   _zz__zz__17_22_inner_macOut_1;
  wire       [15:0]   _zz__17_22_inner_macOut_1;
  wire       [15:0]   _zz__17_22_inner_macOut_2;
  reg        [7:0]    _17_22_inner_activation;
  reg        [7:0]    _17_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_22_inner_macOut;

  assign _zz__zz__17_22_inner_macOut = ($signed(io_mulInput) * $signed(_17_22_inner_activation));
  assign _zz__zz__17_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_22_inner_macOut)) ? 16'h007f : _zz__17_22_inner_macOut_2);
  assign _zz__17_22_inner_macOut_2 = (($signed(_zz__17_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_22_inner_activation;
    end else begin
      io_macOut = _17_22_inner_macOut;
    end
  end

  assign _zz__17_22_inner_macOut = ($signed(_zz__zz__17_22_inner_macOut) + $signed(_zz__zz__17_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_22_inner_activation <= 8'h00;
      _17_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_22_inner_activation <= io_addInput;
      end else begin
        _17_22_inner_macOut <= _zz__17_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_565 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_21_inner_macOut;
  wire       [15:0]   _zz__zz__17_21_inner_macOut_1;
  wire       [15:0]   _zz__17_21_inner_macOut_1;
  wire       [15:0]   _zz__17_21_inner_macOut_2;
  reg        [7:0]    _17_21_inner_activation;
  reg        [7:0]    _17_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_21_inner_macOut;

  assign _zz__zz__17_21_inner_macOut = ($signed(io_mulInput) * $signed(_17_21_inner_activation));
  assign _zz__zz__17_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_21_inner_macOut)) ? 16'h007f : _zz__17_21_inner_macOut_2);
  assign _zz__17_21_inner_macOut_2 = (($signed(_zz__17_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_21_inner_activation;
    end else begin
      io_macOut = _17_21_inner_macOut;
    end
  end

  assign _zz__17_21_inner_macOut = ($signed(_zz__zz__17_21_inner_macOut) + $signed(_zz__zz__17_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_21_inner_activation <= 8'h00;
      _17_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_21_inner_activation <= io_addInput;
      end else begin
        _17_21_inner_macOut <= _zz__17_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_564 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_20_inner_macOut;
  wire       [15:0]   _zz__zz__17_20_inner_macOut_1;
  wire       [15:0]   _zz__17_20_inner_macOut_1;
  wire       [15:0]   _zz__17_20_inner_macOut_2;
  reg        [7:0]    _17_20_inner_activation;
  reg        [7:0]    _17_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_20_inner_macOut;

  assign _zz__zz__17_20_inner_macOut = ($signed(io_mulInput) * $signed(_17_20_inner_activation));
  assign _zz__zz__17_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_20_inner_macOut)) ? 16'h007f : _zz__17_20_inner_macOut_2);
  assign _zz__17_20_inner_macOut_2 = (($signed(_zz__17_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_20_inner_activation;
    end else begin
      io_macOut = _17_20_inner_macOut;
    end
  end

  assign _zz__17_20_inner_macOut = ($signed(_zz__zz__17_20_inner_macOut) + $signed(_zz__zz__17_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_20_inner_activation <= 8'h00;
      _17_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_20_inner_activation <= io_addInput;
      end else begin
        _17_20_inner_macOut <= _zz__17_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_563 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_19_inner_macOut;
  wire       [15:0]   _zz__zz__17_19_inner_macOut_1;
  wire       [15:0]   _zz__17_19_inner_macOut_1;
  wire       [15:0]   _zz__17_19_inner_macOut_2;
  reg        [7:0]    _17_19_inner_activation;
  reg        [7:0]    _17_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_19_inner_macOut;

  assign _zz__zz__17_19_inner_macOut = ($signed(io_mulInput) * $signed(_17_19_inner_activation));
  assign _zz__zz__17_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_19_inner_macOut)) ? 16'h007f : _zz__17_19_inner_macOut_2);
  assign _zz__17_19_inner_macOut_2 = (($signed(_zz__17_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_19_inner_activation;
    end else begin
      io_macOut = _17_19_inner_macOut;
    end
  end

  assign _zz__17_19_inner_macOut = ($signed(_zz__zz__17_19_inner_macOut) + $signed(_zz__zz__17_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_19_inner_activation <= 8'h00;
      _17_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_19_inner_activation <= io_addInput;
      end else begin
        _17_19_inner_macOut <= _zz__17_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_562 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_18_inner_macOut;
  wire       [15:0]   _zz__zz__17_18_inner_macOut_1;
  wire       [15:0]   _zz__17_18_inner_macOut_1;
  wire       [15:0]   _zz__17_18_inner_macOut_2;
  reg        [7:0]    _17_18_inner_activation;
  reg        [7:0]    _17_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_18_inner_macOut;

  assign _zz__zz__17_18_inner_macOut = ($signed(io_mulInput) * $signed(_17_18_inner_activation));
  assign _zz__zz__17_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_18_inner_macOut)) ? 16'h007f : _zz__17_18_inner_macOut_2);
  assign _zz__17_18_inner_macOut_2 = (($signed(_zz__17_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_18_inner_activation;
    end else begin
      io_macOut = _17_18_inner_macOut;
    end
  end

  assign _zz__17_18_inner_macOut = ($signed(_zz__zz__17_18_inner_macOut) + $signed(_zz__zz__17_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_18_inner_activation <= 8'h00;
      _17_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_18_inner_activation <= io_addInput;
      end else begin
        _17_18_inner_macOut <= _zz__17_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_561 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_17_inner_macOut;
  wire       [15:0]   _zz__zz__17_17_inner_macOut_1;
  wire       [15:0]   _zz__17_17_inner_macOut_1;
  wire       [15:0]   _zz__17_17_inner_macOut_2;
  reg        [7:0]    _17_17_inner_activation;
  reg        [7:0]    _17_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_17_inner_macOut;

  assign _zz__zz__17_17_inner_macOut = ($signed(io_mulInput) * $signed(_17_17_inner_activation));
  assign _zz__zz__17_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_17_inner_macOut)) ? 16'h007f : _zz__17_17_inner_macOut_2);
  assign _zz__17_17_inner_macOut_2 = (($signed(_zz__17_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_17_inner_activation;
    end else begin
      io_macOut = _17_17_inner_macOut;
    end
  end

  assign _zz__17_17_inner_macOut = ($signed(_zz__zz__17_17_inner_macOut) + $signed(_zz__zz__17_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_17_inner_activation <= 8'h00;
      _17_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_17_inner_activation <= io_addInput;
      end else begin
        _17_17_inner_macOut <= _zz__17_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_560 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_16_inner_macOut;
  wire       [15:0]   _zz__zz__17_16_inner_macOut_1;
  wire       [15:0]   _zz__17_16_inner_macOut_1;
  wire       [15:0]   _zz__17_16_inner_macOut_2;
  reg        [7:0]    _17_16_inner_activation;
  reg        [7:0]    _17_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_16_inner_macOut;

  assign _zz__zz__17_16_inner_macOut = ($signed(io_mulInput) * $signed(_17_16_inner_activation));
  assign _zz__zz__17_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_16_inner_macOut)) ? 16'h007f : _zz__17_16_inner_macOut_2);
  assign _zz__17_16_inner_macOut_2 = (($signed(_zz__17_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_16_inner_activation;
    end else begin
      io_macOut = _17_16_inner_macOut;
    end
  end

  assign _zz__17_16_inner_macOut = ($signed(_zz__zz__17_16_inner_macOut) + $signed(_zz__zz__17_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_16_inner_activation <= 8'h00;
      _17_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_16_inner_activation <= io_addInput;
      end else begin
        _17_16_inner_macOut <= _zz__17_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_559 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_15_inner_macOut;
  wire       [15:0]   _zz__zz__17_15_inner_macOut_1;
  wire       [15:0]   _zz__17_15_inner_macOut_1;
  wire       [15:0]   _zz__17_15_inner_macOut_2;
  reg        [7:0]    _17_15_inner_activation;
  reg        [7:0]    _17_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_15_inner_macOut;

  assign _zz__zz__17_15_inner_macOut = ($signed(io_mulInput) * $signed(_17_15_inner_activation));
  assign _zz__zz__17_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_15_inner_macOut)) ? 16'h007f : _zz__17_15_inner_macOut_2);
  assign _zz__17_15_inner_macOut_2 = (($signed(_zz__17_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_15_inner_activation;
    end else begin
      io_macOut = _17_15_inner_macOut;
    end
  end

  assign _zz__17_15_inner_macOut = ($signed(_zz__zz__17_15_inner_macOut) + $signed(_zz__zz__17_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_15_inner_activation <= 8'h00;
      _17_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_15_inner_activation <= io_addInput;
      end else begin
        _17_15_inner_macOut <= _zz__17_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_558 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_14_inner_macOut;
  wire       [15:0]   _zz__zz__17_14_inner_macOut_1;
  wire       [15:0]   _zz__17_14_inner_macOut_1;
  wire       [15:0]   _zz__17_14_inner_macOut_2;
  reg        [7:0]    _17_14_inner_activation;
  reg        [7:0]    _17_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_14_inner_macOut;

  assign _zz__zz__17_14_inner_macOut = ($signed(io_mulInput) * $signed(_17_14_inner_activation));
  assign _zz__zz__17_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_14_inner_macOut)) ? 16'h007f : _zz__17_14_inner_macOut_2);
  assign _zz__17_14_inner_macOut_2 = (($signed(_zz__17_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_14_inner_activation;
    end else begin
      io_macOut = _17_14_inner_macOut;
    end
  end

  assign _zz__17_14_inner_macOut = ($signed(_zz__zz__17_14_inner_macOut) + $signed(_zz__zz__17_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_14_inner_activation <= 8'h00;
      _17_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_14_inner_activation <= io_addInput;
      end else begin
        _17_14_inner_macOut <= _zz__17_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_557 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_13_inner_macOut;
  wire       [15:0]   _zz__zz__17_13_inner_macOut_1;
  wire       [15:0]   _zz__17_13_inner_macOut_1;
  wire       [15:0]   _zz__17_13_inner_macOut_2;
  reg        [7:0]    _17_13_inner_activation;
  reg        [7:0]    _17_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_13_inner_macOut;

  assign _zz__zz__17_13_inner_macOut = ($signed(io_mulInput) * $signed(_17_13_inner_activation));
  assign _zz__zz__17_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_13_inner_macOut)) ? 16'h007f : _zz__17_13_inner_macOut_2);
  assign _zz__17_13_inner_macOut_2 = (($signed(_zz__17_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_13_inner_activation;
    end else begin
      io_macOut = _17_13_inner_macOut;
    end
  end

  assign _zz__17_13_inner_macOut = ($signed(_zz__zz__17_13_inner_macOut) + $signed(_zz__zz__17_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_13_inner_activation <= 8'h00;
      _17_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_13_inner_activation <= io_addInput;
      end else begin
        _17_13_inner_macOut <= _zz__17_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_556 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_12_inner_macOut;
  wire       [15:0]   _zz__zz__17_12_inner_macOut_1;
  wire       [15:0]   _zz__17_12_inner_macOut_1;
  wire       [15:0]   _zz__17_12_inner_macOut_2;
  reg        [7:0]    _17_12_inner_activation;
  reg        [7:0]    _17_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_12_inner_macOut;

  assign _zz__zz__17_12_inner_macOut = ($signed(io_mulInput) * $signed(_17_12_inner_activation));
  assign _zz__zz__17_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_12_inner_macOut)) ? 16'h007f : _zz__17_12_inner_macOut_2);
  assign _zz__17_12_inner_macOut_2 = (($signed(_zz__17_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_12_inner_activation;
    end else begin
      io_macOut = _17_12_inner_macOut;
    end
  end

  assign _zz__17_12_inner_macOut = ($signed(_zz__zz__17_12_inner_macOut) + $signed(_zz__zz__17_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_12_inner_activation <= 8'h00;
      _17_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_12_inner_activation <= io_addInput;
      end else begin
        _17_12_inner_macOut <= _zz__17_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_555 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_11_inner_macOut;
  wire       [15:0]   _zz__zz__17_11_inner_macOut_1;
  wire       [15:0]   _zz__17_11_inner_macOut_1;
  wire       [15:0]   _zz__17_11_inner_macOut_2;
  reg        [7:0]    _17_11_inner_activation;
  reg        [7:0]    _17_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_11_inner_macOut;

  assign _zz__zz__17_11_inner_macOut = ($signed(io_mulInput) * $signed(_17_11_inner_activation));
  assign _zz__zz__17_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_11_inner_macOut)) ? 16'h007f : _zz__17_11_inner_macOut_2);
  assign _zz__17_11_inner_macOut_2 = (($signed(_zz__17_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_11_inner_activation;
    end else begin
      io_macOut = _17_11_inner_macOut;
    end
  end

  assign _zz__17_11_inner_macOut = ($signed(_zz__zz__17_11_inner_macOut) + $signed(_zz__zz__17_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_11_inner_activation <= 8'h00;
      _17_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_11_inner_activation <= io_addInput;
      end else begin
        _17_11_inner_macOut <= _zz__17_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_554 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_10_inner_macOut;
  wire       [15:0]   _zz__zz__17_10_inner_macOut_1;
  wire       [15:0]   _zz__17_10_inner_macOut_1;
  wire       [15:0]   _zz__17_10_inner_macOut_2;
  reg        [7:0]    _17_10_inner_activation;
  reg        [7:0]    _17_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_10_inner_macOut;

  assign _zz__zz__17_10_inner_macOut = ($signed(io_mulInput) * $signed(_17_10_inner_activation));
  assign _zz__zz__17_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_10_inner_macOut)) ? 16'h007f : _zz__17_10_inner_macOut_2);
  assign _zz__17_10_inner_macOut_2 = (($signed(_zz__17_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_10_inner_activation;
    end else begin
      io_macOut = _17_10_inner_macOut;
    end
  end

  assign _zz__17_10_inner_macOut = ($signed(_zz__zz__17_10_inner_macOut) + $signed(_zz__zz__17_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_10_inner_activation <= 8'h00;
      _17_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_10_inner_activation <= io_addInput;
      end else begin
        _17_10_inner_macOut <= _zz__17_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_553 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_9_inner_macOut;
  wire       [15:0]   _zz__zz__17_9_inner_macOut_1;
  wire       [15:0]   _zz__17_9_inner_macOut_1;
  wire       [15:0]   _zz__17_9_inner_macOut_2;
  reg        [7:0]    _17_9_inner_activation;
  reg        [7:0]    _17_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_9_inner_macOut;

  assign _zz__zz__17_9_inner_macOut = ($signed(io_mulInput) * $signed(_17_9_inner_activation));
  assign _zz__zz__17_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_9_inner_macOut)) ? 16'h007f : _zz__17_9_inner_macOut_2);
  assign _zz__17_9_inner_macOut_2 = (($signed(_zz__17_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_9_inner_activation;
    end else begin
      io_macOut = _17_9_inner_macOut;
    end
  end

  assign _zz__17_9_inner_macOut = ($signed(_zz__zz__17_9_inner_macOut) + $signed(_zz__zz__17_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_9_inner_activation <= 8'h00;
      _17_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_9_inner_activation <= io_addInput;
      end else begin
        _17_9_inner_macOut <= _zz__17_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_552 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_8_inner_macOut;
  wire       [15:0]   _zz__zz__17_8_inner_macOut_1;
  wire       [15:0]   _zz__17_8_inner_macOut_1;
  wire       [15:0]   _zz__17_8_inner_macOut_2;
  reg        [7:0]    _17_8_inner_activation;
  reg        [7:0]    _17_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_8_inner_macOut;

  assign _zz__zz__17_8_inner_macOut = ($signed(io_mulInput) * $signed(_17_8_inner_activation));
  assign _zz__zz__17_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_8_inner_macOut)) ? 16'h007f : _zz__17_8_inner_macOut_2);
  assign _zz__17_8_inner_macOut_2 = (($signed(_zz__17_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_8_inner_activation;
    end else begin
      io_macOut = _17_8_inner_macOut;
    end
  end

  assign _zz__17_8_inner_macOut = ($signed(_zz__zz__17_8_inner_macOut) + $signed(_zz__zz__17_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_8_inner_activation <= 8'h00;
      _17_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_8_inner_activation <= io_addInput;
      end else begin
        _17_8_inner_macOut <= _zz__17_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_551 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_7_inner_macOut;
  wire       [15:0]   _zz__zz__17_7_inner_macOut_1;
  wire       [15:0]   _zz__17_7_inner_macOut_1;
  wire       [15:0]   _zz__17_7_inner_macOut_2;
  reg        [7:0]    _17_7_inner_activation;
  reg        [7:0]    _17_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_7_inner_macOut;

  assign _zz__zz__17_7_inner_macOut = ($signed(io_mulInput) * $signed(_17_7_inner_activation));
  assign _zz__zz__17_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_7_inner_macOut)) ? 16'h007f : _zz__17_7_inner_macOut_2);
  assign _zz__17_7_inner_macOut_2 = (($signed(_zz__17_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_7_inner_activation;
    end else begin
      io_macOut = _17_7_inner_macOut;
    end
  end

  assign _zz__17_7_inner_macOut = ($signed(_zz__zz__17_7_inner_macOut) + $signed(_zz__zz__17_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_7_inner_activation <= 8'h00;
      _17_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_7_inner_activation <= io_addInput;
      end else begin
        _17_7_inner_macOut <= _zz__17_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_550 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_6_inner_macOut;
  wire       [15:0]   _zz__zz__17_6_inner_macOut_1;
  wire       [15:0]   _zz__17_6_inner_macOut_1;
  wire       [15:0]   _zz__17_6_inner_macOut_2;
  reg        [7:0]    _17_6_inner_activation;
  reg        [7:0]    _17_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_6_inner_macOut;

  assign _zz__zz__17_6_inner_macOut = ($signed(io_mulInput) * $signed(_17_6_inner_activation));
  assign _zz__zz__17_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_6_inner_macOut)) ? 16'h007f : _zz__17_6_inner_macOut_2);
  assign _zz__17_6_inner_macOut_2 = (($signed(_zz__17_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_6_inner_activation;
    end else begin
      io_macOut = _17_6_inner_macOut;
    end
  end

  assign _zz__17_6_inner_macOut = ($signed(_zz__zz__17_6_inner_macOut) + $signed(_zz__zz__17_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_6_inner_activation <= 8'h00;
      _17_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_6_inner_activation <= io_addInput;
      end else begin
        _17_6_inner_macOut <= _zz__17_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_549 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_5_inner_macOut;
  wire       [15:0]   _zz__zz__17_5_inner_macOut_1;
  wire       [15:0]   _zz__17_5_inner_macOut_1;
  wire       [15:0]   _zz__17_5_inner_macOut_2;
  reg        [7:0]    _17_5_inner_activation;
  reg        [7:0]    _17_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_5_inner_macOut;

  assign _zz__zz__17_5_inner_macOut = ($signed(io_mulInput) * $signed(_17_5_inner_activation));
  assign _zz__zz__17_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_5_inner_macOut)) ? 16'h007f : _zz__17_5_inner_macOut_2);
  assign _zz__17_5_inner_macOut_2 = (($signed(_zz__17_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_5_inner_activation;
    end else begin
      io_macOut = _17_5_inner_macOut;
    end
  end

  assign _zz__17_5_inner_macOut = ($signed(_zz__zz__17_5_inner_macOut) + $signed(_zz__zz__17_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_5_inner_activation <= 8'h00;
      _17_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_5_inner_activation <= io_addInput;
      end else begin
        _17_5_inner_macOut <= _zz__17_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_548 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_4_inner_macOut;
  wire       [15:0]   _zz__zz__17_4_inner_macOut_1;
  wire       [15:0]   _zz__17_4_inner_macOut_1;
  wire       [15:0]   _zz__17_4_inner_macOut_2;
  reg        [7:0]    _17_4_inner_activation;
  reg        [7:0]    _17_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_4_inner_macOut;

  assign _zz__zz__17_4_inner_macOut = ($signed(io_mulInput) * $signed(_17_4_inner_activation));
  assign _zz__zz__17_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_4_inner_macOut)) ? 16'h007f : _zz__17_4_inner_macOut_2);
  assign _zz__17_4_inner_macOut_2 = (($signed(_zz__17_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_4_inner_activation;
    end else begin
      io_macOut = _17_4_inner_macOut;
    end
  end

  assign _zz__17_4_inner_macOut = ($signed(_zz__zz__17_4_inner_macOut) + $signed(_zz__zz__17_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_4_inner_activation <= 8'h00;
      _17_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_4_inner_activation <= io_addInput;
      end else begin
        _17_4_inner_macOut <= _zz__17_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_547 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_3_inner_macOut;
  wire       [15:0]   _zz__zz__17_3_inner_macOut_1;
  wire       [15:0]   _zz__17_3_inner_macOut_1;
  wire       [15:0]   _zz__17_3_inner_macOut_2;
  reg        [7:0]    _17_3_inner_activation;
  reg        [7:0]    _17_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_3_inner_macOut;

  assign _zz__zz__17_3_inner_macOut = ($signed(io_mulInput) * $signed(_17_3_inner_activation));
  assign _zz__zz__17_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_3_inner_macOut)) ? 16'h007f : _zz__17_3_inner_macOut_2);
  assign _zz__17_3_inner_macOut_2 = (($signed(_zz__17_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_3_inner_activation;
    end else begin
      io_macOut = _17_3_inner_macOut;
    end
  end

  assign _zz__17_3_inner_macOut = ($signed(_zz__zz__17_3_inner_macOut) + $signed(_zz__zz__17_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_3_inner_activation <= 8'h00;
      _17_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_3_inner_activation <= io_addInput;
      end else begin
        _17_3_inner_macOut <= _zz__17_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_546 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_2_inner_macOut;
  wire       [15:0]   _zz__zz__17_2_inner_macOut_1;
  wire       [15:0]   _zz__17_2_inner_macOut_1;
  wire       [15:0]   _zz__17_2_inner_macOut_2;
  reg        [7:0]    _17_2_inner_activation;
  reg        [7:0]    _17_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_2_inner_macOut;

  assign _zz__zz__17_2_inner_macOut = ($signed(io_mulInput) * $signed(_17_2_inner_activation));
  assign _zz__zz__17_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_2_inner_macOut)) ? 16'h007f : _zz__17_2_inner_macOut_2);
  assign _zz__17_2_inner_macOut_2 = (($signed(_zz__17_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_2_inner_activation;
    end else begin
      io_macOut = _17_2_inner_macOut;
    end
  end

  assign _zz__17_2_inner_macOut = ($signed(_zz__zz__17_2_inner_macOut) + $signed(_zz__zz__17_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_2_inner_activation <= 8'h00;
      _17_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_2_inner_activation <= io_addInput;
      end else begin
        _17_2_inner_macOut <= _zz__17_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_545 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_1_inner_macOut;
  wire       [15:0]   _zz__zz__17_1_inner_macOut_1;
  wire       [15:0]   _zz__17_1_inner_macOut_1;
  wire       [15:0]   _zz__17_1_inner_macOut_2;
  reg        [7:0]    _17_1_inner_activation;
  reg        [7:0]    _17_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_1_inner_macOut;

  assign _zz__zz__17_1_inner_macOut = ($signed(io_mulInput) * $signed(_17_1_inner_activation));
  assign _zz__zz__17_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_1_inner_macOut)) ? 16'h007f : _zz__17_1_inner_macOut_2);
  assign _zz__17_1_inner_macOut_2 = (($signed(_zz__17_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_1_inner_activation;
    end else begin
      io_macOut = _17_1_inner_macOut;
    end
  end

  assign _zz__17_1_inner_macOut = ($signed(_zz__zz__17_1_inner_macOut) + $signed(_zz__zz__17_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_1_inner_activation <= 8'h00;
      _17_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_1_inner_activation <= io_addInput;
      end else begin
        _17_1_inner_macOut <= _zz__17_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_544 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__17_0_inner_macOut;
  wire       [15:0]   _zz__zz__17_0_inner_macOut_1;
  wire       [15:0]   _zz__17_0_inner_macOut_1;
  wire       [15:0]   _zz__17_0_inner_macOut_2;
  reg        [7:0]    _17_0_inner_activation;
  reg        [7:0]    _17_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__17_0_inner_macOut;

  assign _zz__zz__17_0_inner_macOut = ($signed(io_mulInput) * $signed(_17_0_inner_activation));
  assign _zz__zz__17_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__17_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__17_0_inner_macOut)) ? 16'h007f : _zz__17_0_inner_macOut_2);
  assign _zz__17_0_inner_macOut_2 = (($signed(_zz__17_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__17_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _17_0_inner_activation;
    end else begin
      io_macOut = _17_0_inner_macOut;
    end
  end

  assign _zz__17_0_inner_macOut = ($signed(_zz__zz__17_0_inner_macOut) + $signed(_zz__zz__17_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _17_0_inner_activation <= 8'h00;
      _17_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _17_0_inner_activation <= io_addInput;
      end else begin
        _17_0_inner_macOut <= _zz__17_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_543 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_31_inner_macOut;
  wire       [15:0]   _zz__zz__16_31_inner_macOut_1;
  wire       [15:0]   _zz__16_31_inner_macOut_1;
  wire       [15:0]   _zz__16_31_inner_macOut_2;
  reg        [7:0]    _16_31_inner_activation;
  reg        [7:0]    _16_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_31_inner_macOut;

  assign _zz__zz__16_31_inner_macOut = ($signed(io_mulInput) * $signed(_16_31_inner_activation));
  assign _zz__zz__16_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_31_inner_macOut)) ? 16'h007f : _zz__16_31_inner_macOut_2);
  assign _zz__16_31_inner_macOut_2 = (($signed(_zz__16_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_31_inner_activation;
    end else begin
      io_macOut = _16_31_inner_macOut;
    end
  end

  assign _zz__16_31_inner_macOut = ($signed(_zz__zz__16_31_inner_macOut) + $signed(_zz__zz__16_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_31_inner_activation <= 8'h00;
      _16_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_31_inner_activation <= io_addInput;
      end else begin
        _16_31_inner_macOut <= _zz__16_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_542 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_30_inner_macOut;
  wire       [15:0]   _zz__zz__16_30_inner_macOut_1;
  wire       [15:0]   _zz__16_30_inner_macOut_1;
  wire       [15:0]   _zz__16_30_inner_macOut_2;
  reg        [7:0]    _16_30_inner_activation;
  reg        [7:0]    _16_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_30_inner_macOut;

  assign _zz__zz__16_30_inner_macOut = ($signed(io_mulInput) * $signed(_16_30_inner_activation));
  assign _zz__zz__16_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_30_inner_macOut)) ? 16'h007f : _zz__16_30_inner_macOut_2);
  assign _zz__16_30_inner_macOut_2 = (($signed(_zz__16_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_30_inner_activation;
    end else begin
      io_macOut = _16_30_inner_macOut;
    end
  end

  assign _zz__16_30_inner_macOut = ($signed(_zz__zz__16_30_inner_macOut) + $signed(_zz__zz__16_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_30_inner_activation <= 8'h00;
      _16_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_30_inner_activation <= io_addInput;
      end else begin
        _16_30_inner_macOut <= _zz__16_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_541 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_29_inner_macOut;
  wire       [15:0]   _zz__zz__16_29_inner_macOut_1;
  wire       [15:0]   _zz__16_29_inner_macOut_1;
  wire       [15:0]   _zz__16_29_inner_macOut_2;
  reg        [7:0]    _16_29_inner_activation;
  reg        [7:0]    _16_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_29_inner_macOut;

  assign _zz__zz__16_29_inner_macOut = ($signed(io_mulInput) * $signed(_16_29_inner_activation));
  assign _zz__zz__16_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_29_inner_macOut)) ? 16'h007f : _zz__16_29_inner_macOut_2);
  assign _zz__16_29_inner_macOut_2 = (($signed(_zz__16_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_29_inner_activation;
    end else begin
      io_macOut = _16_29_inner_macOut;
    end
  end

  assign _zz__16_29_inner_macOut = ($signed(_zz__zz__16_29_inner_macOut) + $signed(_zz__zz__16_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_29_inner_activation <= 8'h00;
      _16_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_29_inner_activation <= io_addInput;
      end else begin
        _16_29_inner_macOut <= _zz__16_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_540 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_28_inner_macOut;
  wire       [15:0]   _zz__zz__16_28_inner_macOut_1;
  wire       [15:0]   _zz__16_28_inner_macOut_1;
  wire       [15:0]   _zz__16_28_inner_macOut_2;
  reg        [7:0]    _16_28_inner_activation;
  reg        [7:0]    _16_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_28_inner_macOut;

  assign _zz__zz__16_28_inner_macOut = ($signed(io_mulInput) * $signed(_16_28_inner_activation));
  assign _zz__zz__16_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_28_inner_macOut)) ? 16'h007f : _zz__16_28_inner_macOut_2);
  assign _zz__16_28_inner_macOut_2 = (($signed(_zz__16_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_28_inner_activation;
    end else begin
      io_macOut = _16_28_inner_macOut;
    end
  end

  assign _zz__16_28_inner_macOut = ($signed(_zz__zz__16_28_inner_macOut) + $signed(_zz__zz__16_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_28_inner_activation <= 8'h00;
      _16_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_28_inner_activation <= io_addInput;
      end else begin
        _16_28_inner_macOut <= _zz__16_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_539 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_27_inner_macOut;
  wire       [15:0]   _zz__zz__16_27_inner_macOut_1;
  wire       [15:0]   _zz__16_27_inner_macOut_1;
  wire       [15:0]   _zz__16_27_inner_macOut_2;
  reg        [7:0]    _16_27_inner_activation;
  reg        [7:0]    _16_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_27_inner_macOut;

  assign _zz__zz__16_27_inner_macOut = ($signed(io_mulInput) * $signed(_16_27_inner_activation));
  assign _zz__zz__16_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_27_inner_macOut)) ? 16'h007f : _zz__16_27_inner_macOut_2);
  assign _zz__16_27_inner_macOut_2 = (($signed(_zz__16_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_27_inner_activation;
    end else begin
      io_macOut = _16_27_inner_macOut;
    end
  end

  assign _zz__16_27_inner_macOut = ($signed(_zz__zz__16_27_inner_macOut) + $signed(_zz__zz__16_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_27_inner_activation <= 8'h00;
      _16_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_27_inner_activation <= io_addInput;
      end else begin
        _16_27_inner_macOut <= _zz__16_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_538 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_26_inner_macOut;
  wire       [15:0]   _zz__zz__16_26_inner_macOut_1;
  wire       [15:0]   _zz__16_26_inner_macOut_1;
  wire       [15:0]   _zz__16_26_inner_macOut_2;
  reg        [7:0]    _16_26_inner_activation;
  reg        [7:0]    _16_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_26_inner_macOut;

  assign _zz__zz__16_26_inner_macOut = ($signed(io_mulInput) * $signed(_16_26_inner_activation));
  assign _zz__zz__16_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_26_inner_macOut)) ? 16'h007f : _zz__16_26_inner_macOut_2);
  assign _zz__16_26_inner_macOut_2 = (($signed(_zz__16_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_26_inner_activation;
    end else begin
      io_macOut = _16_26_inner_macOut;
    end
  end

  assign _zz__16_26_inner_macOut = ($signed(_zz__zz__16_26_inner_macOut) + $signed(_zz__zz__16_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_26_inner_activation <= 8'h00;
      _16_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_26_inner_activation <= io_addInput;
      end else begin
        _16_26_inner_macOut <= _zz__16_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_537 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_25_inner_macOut;
  wire       [15:0]   _zz__zz__16_25_inner_macOut_1;
  wire       [15:0]   _zz__16_25_inner_macOut_1;
  wire       [15:0]   _zz__16_25_inner_macOut_2;
  reg        [7:0]    _16_25_inner_activation;
  reg        [7:0]    _16_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_25_inner_macOut;

  assign _zz__zz__16_25_inner_macOut = ($signed(io_mulInput) * $signed(_16_25_inner_activation));
  assign _zz__zz__16_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_25_inner_macOut)) ? 16'h007f : _zz__16_25_inner_macOut_2);
  assign _zz__16_25_inner_macOut_2 = (($signed(_zz__16_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_25_inner_activation;
    end else begin
      io_macOut = _16_25_inner_macOut;
    end
  end

  assign _zz__16_25_inner_macOut = ($signed(_zz__zz__16_25_inner_macOut) + $signed(_zz__zz__16_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_25_inner_activation <= 8'h00;
      _16_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_25_inner_activation <= io_addInput;
      end else begin
        _16_25_inner_macOut <= _zz__16_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_536 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_24_inner_macOut;
  wire       [15:0]   _zz__zz__16_24_inner_macOut_1;
  wire       [15:0]   _zz__16_24_inner_macOut_1;
  wire       [15:0]   _zz__16_24_inner_macOut_2;
  reg        [7:0]    _16_24_inner_activation;
  reg        [7:0]    _16_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_24_inner_macOut;

  assign _zz__zz__16_24_inner_macOut = ($signed(io_mulInput) * $signed(_16_24_inner_activation));
  assign _zz__zz__16_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_24_inner_macOut)) ? 16'h007f : _zz__16_24_inner_macOut_2);
  assign _zz__16_24_inner_macOut_2 = (($signed(_zz__16_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_24_inner_activation;
    end else begin
      io_macOut = _16_24_inner_macOut;
    end
  end

  assign _zz__16_24_inner_macOut = ($signed(_zz__zz__16_24_inner_macOut) + $signed(_zz__zz__16_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_24_inner_activation <= 8'h00;
      _16_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_24_inner_activation <= io_addInput;
      end else begin
        _16_24_inner_macOut <= _zz__16_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_535 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_23_inner_macOut;
  wire       [15:0]   _zz__zz__16_23_inner_macOut_1;
  wire       [15:0]   _zz__16_23_inner_macOut_1;
  wire       [15:0]   _zz__16_23_inner_macOut_2;
  reg        [7:0]    _16_23_inner_activation;
  reg        [7:0]    _16_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_23_inner_macOut;

  assign _zz__zz__16_23_inner_macOut = ($signed(io_mulInput) * $signed(_16_23_inner_activation));
  assign _zz__zz__16_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_23_inner_macOut)) ? 16'h007f : _zz__16_23_inner_macOut_2);
  assign _zz__16_23_inner_macOut_2 = (($signed(_zz__16_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_23_inner_activation;
    end else begin
      io_macOut = _16_23_inner_macOut;
    end
  end

  assign _zz__16_23_inner_macOut = ($signed(_zz__zz__16_23_inner_macOut) + $signed(_zz__zz__16_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_23_inner_activation <= 8'h00;
      _16_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_23_inner_activation <= io_addInput;
      end else begin
        _16_23_inner_macOut <= _zz__16_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_534 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_22_inner_macOut;
  wire       [15:0]   _zz__zz__16_22_inner_macOut_1;
  wire       [15:0]   _zz__16_22_inner_macOut_1;
  wire       [15:0]   _zz__16_22_inner_macOut_2;
  reg        [7:0]    _16_22_inner_activation;
  reg        [7:0]    _16_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_22_inner_macOut;

  assign _zz__zz__16_22_inner_macOut = ($signed(io_mulInput) * $signed(_16_22_inner_activation));
  assign _zz__zz__16_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_22_inner_macOut)) ? 16'h007f : _zz__16_22_inner_macOut_2);
  assign _zz__16_22_inner_macOut_2 = (($signed(_zz__16_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_22_inner_activation;
    end else begin
      io_macOut = _16_22_inner_macOut;
    end
  end

  assign _zz__16_22_inner_macOut = ($signed(_zz__zz__16_22_inner_macOut) + $signed(_zz__zz__16_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_22_inner_activation <= 8'h00;
      _16_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_22_inner_activation <= io_addInput;
      end else begin
        _16_22_inner_macOut <= _zz__16_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_533 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_21_inner_macOut;
  wire       [15:0]   _zz__zz__16_21_inner_macOut_1;
  wire       [15:0]   _zz__16_21_inner_macOut_1;
  wire       [15:0]   _zz__16_21_inner_macOut_2;
  reg        [7:0]    _16_21_inner_activation;
  reg        [7:0]    _16_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_21_inner_macOut;

  assign _zz__zz__16_21_inner_macOut = ($signed(io_mulInput) * $signed(_16_21_inner_activation));
  assign _zz__zz__16_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_21_inner_macOut)) ? 16'h007f : _zz__16_21_inner_macOut_2);
  assign _zz__16_21_inner_macOut_2 = (($signed(_zz__16_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_21_inner_activation;
    end else begin
      io_macOut = _16_21_inner_macOut;
    end
  end

  assign _zz__16_21_inner_macOut = ($signed(_zz__zz__16_21_inner_macOut) + $signed(_zz__zz__16_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_21_inner_activation <= 8'h00;
      _16_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_21_inner_activation <= io_addInput;
      end else begin
        _16_21_inner_macOut <= _zz__16_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_532 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_20_inner_macOut;
  wire       [15:0]   _zz__zz__16_20_inner_macOut_1;
  wire       [15:0]   _zz__16_20_inner_macOut_1;
  wire       [15:0]   _zz__16_20_inner_macOut_2;
  reg        [7:0]    _16_20_inner_activation;
  reg        [7:0]    _16_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_20_inner_macOut;

  assign _zz__zz__16_20_inner_macOut = ($signed(io_mulInput) * $signed(_16_20_inner_activation));
  assign _zz__zz__16_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_20_inner_macOut)) ? 16'h007f : _zz__16_20_inner_macOut_2);
  assign _zz__16_20_inner_macOut_2 = (($signed(_zz__16_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_20_inner_activation;
    end else begin
      io_macOut = _16_20_inner_macOut;
    end
  end

  assign _zz__16_20_inner_macOut = ($signed(_zz__zz__16_20_inner_macOut) + $signed(_zz__zz__16_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_20_inner_activation <= 8'h00;
      _16_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_20_inner_activation <= io_addInput;
      end else begin
        _16_20_inner_macOut <= _zz__16_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_531 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_19_inner_macOut;
  wire       [15:0]   _zz__zz__16_19_inner_macOut_1;
  wire       [15:0]   _zz__16_19_inner_macOut_1;
  wire       [15:0]   _zz__16_19_inner_macOut_2;
  reg        [7:0]    _16_19_inner_activation;
  reg        [7:0]    _16_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_19_inner_macOut;

  assign _zz__zz__16_19_inner_macOut = ($signed(io_mulInput) * $signed(_16_19_inner_activation));
  assign _zz__zz__16_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_19_inner_macOut)) ? 16'h007f : _zz__16_19_inner_macOut_2);
  assign _zz__16_19_inner_macOut_2 = (($signed(_zz__16_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_19_inner_activation;
    end else begin
      io_macOut = _16_19_inner_macOut;
    end
  end

  assign _zz__16_19_inner_macOut = ($signed(_zz__zz__16_19_inner_macOut) + $signed(_zz__zz__16_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_19_inner_activation <= 8'h00;
      _16_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_19_inner_activation <= io_addInput;
      end else begin
        _16_19_inner_macOut <= _zz__16_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_530 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_18_inner_macOut;
  wire       [15:0]   _zz__zz__16_18_inner_macOut_1;
  wire       [15:0]   _zz__16_18_inner_macOut_1;
  wire       [15:0]   _zz__16_18_inner_macOut_2;
  reg        [7:0]    _16_18_inner_activation;
  reg        [7:0]    _16_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_18_inner_macOut;

  assign _zz__zz__16_18_inner_macOut = ($signed(io_mulInput) * $signed(_16_18_inner_activation));
  assign _zz__zz__16_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_18_inner_macOut)) ? 16'h007f : _zz__16_18_inner_macOut_2);
  assign _zz__16_18_inner_macOut_2 = (($signed(_zz__16_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_18_inner_activation;
    end else begin
      io_macOut = _16_18_inner_macOut;
    end
  end

  assign _zz__16_18_inner_macOut = ($signed(_zz__zz__16_18_inner_macOut) + $signed(_zz__zz__16_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_18_inner_activation <= 8'h00;
      _16_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_18_inner_activation <= io_addInput;
      end else begin
        _16_18_inner_macOut <= _zz__16_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_529 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_17_inner_macOut;
  wire       [15:0]   _zz__zz__16_17_inner_macOut_1;
  wire       [15:0]   _zz__16_17_inner_macOut_1;
  wire       [15:0]   _zz__16_17_inner_macOut_2;
  reg        [7:0]    _16_17_inner_activation;
  reg        [7:0]    _16_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_17_inner_macOut;

  assign _zz__zz__16_17_inner_macOut = ($signed(io_mulInput) * $signed(_16_17_inner_activation));
  assign _zz__zz__16_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_17_inner_macOut)) ? 16'h007f : _zz__16_17_inner_macOut_2);
  assign _zz__16_17_inner_macOut_2 = (($signed(_zz__16_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_17_inner_activation;
    end else begin
      io_macOut = _16_17_inner_macOut;
    end
  end

  assign _zz__16_17_inner_macOut = ($signed(_zz__zz__16_17_inner_macOut) + $signed(_zz__zz__16_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_17_inner_activation <= 8'h00;
      _16_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_17_inner_activation <= io_addInput;
      end else begin
        _16_17_inner_macOut <= _zz__16_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_528 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_16_inner_macOut;
  wire       [15:0]   _zz__zz__16_16_inner_macOut_1;
  wire       [15:0]   _zz__16_16_inner_macOut_1;
  wire       [15:0]   _zz__16_16_inner_macOut_2;
  reg        [7:0]    _16_16_inner_activation;
  reg        [7:0]    _16_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_16_inner_macOut;

  assign _zz__zz__16_16_inner_macOut = ($signed(io_mulInput) * $signed(_16_16_inner_activation));
  assign _zz__zz__16_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_16_inner_macOut)) ? 16'h007f : _zz__16_16_inner_macOut_2);
  assign _zz__16_16_inner_macOut_2 = (($signed(_zz__16_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_16_inner_activation;
    end else begin
      io_macOut = _16_16_inner_macOut;
    end
  end

  assign _zz__16_16_inner_macOut = ($signed(_zz__zz__16_16_inner_macOut) + $signed(_zz__zz__16_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_16_inner_activation <= 8'h00;
      _16_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_16_inner_activation <= io_addInput;
      end else begin
        _16_16_inner_macOut <= _zz__16_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_527 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_15_inner_macOut;
  wire       [15:0]   _zz__zz__16_15_inner_macOut_1;
  wire       [15:0]   _zz__16_15_inner_macOut_1;
  wire       [15:0]   _zz__16_15_inner_macOut_2;
  reg        [7:0]    _16_15_inner_activation;
  reg        [7:0]    _16_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_15_inner_macOut;

  assign _zz__zz__16_15_inner_macOut = ($signed(io_mulInput) * $signed(_16_15_inner_activation));
  assign _zz__zz__16_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_15_inner_macOut)) ? 16'h007f : _zz__16_15_inner_macOut_2);
  assign _zz__16_15_inner_macOut_2 = (($signed(_zz__16_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_15_inner_activation;
    end else begin
      io_macOut = _16_15_inner_macOut;
    end
  end

  assign _zz__16_15_inner_macOut = ($signed(_zz__zz__16_15_inner_macOut) + $signed(_zz__zz__16_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_15_inner_activation <= 8'h00;
      _16_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_15_inner_activation <= io_addInput;
      end else begin
        _16_15_inner_macOut <= _zz__16_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_526 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_14_inner_macOut;
  wire       [15:0]   _zz__zz__16_14_inner_macOut_1;
  wire       [15:0]   _zz__16_14_inner_macOut_1;
  wire       [15:0]   _zz__16_14_inner_macOut_2;
  reg        [7:0]    _16_14_inner_activation;
  reg        [7:0]    _16_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_14_inner_macOut;

  assign _zz__zz__16_14_inner_macOut = ($signed(io_mulInput) * $signed(_16_14_inner_activation));
  assign _zz__zz__16_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_14_inner_macOut)) ? 16'h007f : _zz__16_14_inner_macOut_2);
  assign _zz__16_14_inner_macOut_2 = (($signed(_zz__16_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_14_inner_activation;
    end else begin
      io_macOut = _16_14_inner_macOut;
    end
  end

  assign _zz__16_14_inner_macOut = ($signed(_zz__zz__16_14_inner_macOut) + $signed(_zz__zz__16_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_14_inner_activation <= 8'h00;
      _16_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_14_inner_activation <= io_addInput;
      end else begin
        _16_14_inner_macOut <= _zz__16_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_525 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_13_inner_macOut;
  wire       [15:0]   _zz__zz__16_13_inner_macOut_1;
  wire       [15:0]   _zz__16_13_inner_macOut_1;
  wire       [15:0]   _zz__16_13_inner_macOut_2;
  reg        [7:0]    _16_13_inner_activation;
  reg        [7:0]    _16_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_13_inner_macOut;

  assign _zz__zz__16_13_inner_macOut = ($signed(io_mulInput) * $signed(_16_13_inner_activation));
  assign _zz__zz__16_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_13_inner_macOut)) ? 16'h007f : _zz__16_13_inner_macOut_2);
  assign _zz__16_13_inner_macOut_2 = (($signed(_zz__16_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_13_inner_activation;
    end else begin
      io_macOut = _16_13_inner_macOut;
    end
  end

  assign _zz__16_13_inner_macOut = ($signed(_zz__zz__16_13_inner_macOut) + $signed(_zz__zz__16_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_13_inner_activation <= 8'h00;
      _16_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_13_inner_activation <= io_addInput;
      end else begin
        _16_13_inner_macOut <= _zz__16_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_524 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_12_inner_macOut;
  wire       [15:0]   _zz__zz__16_12_inner_macOut_1;
  wire       [15:0]   _zz__16_12_inner_macOut_1;
  wire       [15:0]   _zz__16_12_inner_macOut_2;
  reg        [7:0]    _16_12_inner_activation;
  reg        [7:0]    _16_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_12_inner_macOut;

  assign _zz__zz__16_12_inner_macOut = ($signed(io_mulInput) * $signed(_16_12_inner_activation));
  assign _zz__zz__16_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_12_inner_macOut)) ? 16'h007f : _zz__16_12_inner_macOut_2);
  assign _zz__16_12_inner_macOut_2 = (($signed(_zz__16_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_12_inner_activation;
    end else begin
      io_macOut = _16_12_inner_macOut;
    end
  end

  assign _zz__16_12_inner_macOut = ($signed(_zz__zz__16_12_inner_macOut) + $signed(_zz__zz__16_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_12_inner_activation <= 8'h00;
      _16_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_12_inner_activation <= io_addInput;
      end else begin
        _16_12_inner_macOut <= _zz__16_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_523 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_11_inner_macOut;
  wire       [15:0]   _zz__zz__16_11_inner_macOut_1;
  wire       [15:0]   _zz__16_11_inner_macOut_1;
  wire       [15:0]   _zz__16_11_inner_macOut_2;
  reg        [7:0]    _16_11_inner_activation;
  reg        [7:0]    _16_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_11_inner_macOut;

  assign _zz__zz__16_11_inner_macOut = ($signed(io_mulInput) * $signed(_16_11_inner_activation));
  assign _zz__zz__16_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_11_inner_macOut)) ? 16'h007f : _zz__16_11_inner_macOut_2);
  assign _zz__16_11_inner_macOut_2 = (($signed(_zz__16_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_11_inner_activation;
    end else begin
      io_macOut = _16_11_inner_macOut;
    end
  end

  assign _zz__16_11_inner_macOut = ($signed(_zz__zz__16_11_inner_macOut) + $signed(_zz__zz__16_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_11_inner_activation <= 8'h00;
      _16_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_11_inner_activation <= io_addInput;
      end else begin
        _16_11_inner_macOut <= _zz__16_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_522 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_10_inner_macOut;
  wire       [15:0]   _zz__zz__16_10_inner_macOut_1;
  wire       [15:0]   _zz__16_10_inner_macOut_1;
  wire       [15:0]   _zz__16_10_inner_macOut_2;
  reg        [7:0]    _16_10_inner_activation;
  reg        [7:0]    _16_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_10_inner_macOut;

  assign _zz__zz__16_10_inner_macOut = ($signed(io_mulInput) * $signed(_16_10_inner_activation));
  assign _zz__zz__16_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_10_inner_macOut)) ? 16'h007f : _zz__16_10_inner_macOut_2);
  assign _zz__16_10_inner_macOut_2 = (($signed(_zz__16_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_10_inner_activation;
    end else begin
      io_macOut = _16_10_inner_macOut;
    end
  end

  assign _zz__16_10_inner_macOut = ($signed(_zz__zz__16_10_inner_macOut) + $signed(_zz__zz__16_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_10_inner_activation <= 8'h00;
      _16_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_10_inner_activation <= io_addInput;
      end else begin
        _16_10_inner_macOut <= _zz__16_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_521 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_9_inner_macOut;
  wire       [15:0]   _zz__zz__16_9_inner_macOut_1;
  wire       [15:0]   _zz__16_9_inner_macOut_1;
  wire       [15:0]   _zz__16_9_inner_macOut_2;
  reg        [7:0]    _16_9_inner_activation;
  reg        [7:0]    _16_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_9_inner_macOut;

  assign _zz__zz__16_9_inner_macOut = ($signed(io_mulInput) * $signed(_16_9_inner_activation));
  assign _zz__zz__16_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_9_inner_macOut)) ? 16'h007f : _zz__16_9_inner_macOut_2);
  assign _zz__16_9_inner_macOut_2 = (($signed(_zz__16_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_9_inner_activation;
    end else begin
      io_macOut = _16_9_inner_macOut;
    end
  end

  assign _zz__16_9_inner_macOut = ($signed(_zz__zz__16_9_inner_macOut) + $signed(_zz__zz__16_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_9_inner_activation <= 8'h00;
      _16_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_9_inner_activation <= io_addInput;
      end else begin
        _16_9_inner_macOut <= _zz__16_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_520 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_8_inner_macOut;
  wire       [15:0]   _zz__zz__16_8_inner_macOut_1;
  wire       [15:0]   _zz__16_8_inner_macOut_1;
  wire       [15:0]   _zz__16_8_inner_macOut_2;
  reg        [7:0]    _16_8_inner_activation;
  reg        [7:0]    _16_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_8_inner_macOut;

  assign _zz__zz__16_8_inner_macOut = ($signed(io_mulInput) * $signed(_16_8_inner_activation));
  assign _zz__zz__16_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_8_inner_macOut)) ? 16'h007f : _zz__16_8_inner_macOut_2);
  assign _zz__16_8_inner_macOut_2 = (($signed(_zz__16_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_8_inner_activation;
    end else begin
      io_macOut = _16_8_inner_macOut;
    end
  end

  assign _zz__16_8_inner_macOut = ($signed(_zz__zz__16_8_inner_macOut) + $signed(_zz__zz__16_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_8_inner_activation <= 8'h00;
      _16_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_8_inner_activation <= io_addInput;
      end else begin
        _16_8_inner_macOut <= _zz__16_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_519 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_7_inner_macOut;
  wire       [15:0]   _zz__zz__16_7_inner_macOut_1;
  wire       [15:0]   _zz__16_7_inner_macOut_1;
  wire       [15:0]   _zz__16_7_inner_macOut_2;
  reg        [7:0]    _16_7_inner_activation;
  reg        [7:0]    _16_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_7_inner_macOut;

  assign _zz__zz__16_7_inner_macOut = ($signed(io_mulInput) * $signed(_16_7_inner_activation));
  assign _zz__zz__16_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_7_inner_macOut)) ? 16'h007f : _zz__16_7_inner_macOut_2);
  assign _zz__16_7_inner_macOut_2 = (($signed(_zz__16_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_7_inner_activation;
    end else begin
      io_macOut = _16_7_inner_macOut;
    end
  end

  assign _zz__16_7_inner_macOut = ($signed(_zz__zz__16_7_inner_macOut) + $signed(_zz__zz__16_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_7_inner_activation <= 8'h00;
      _16_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_7_inner_activation <= io_addInput;
      end else begin
        _16_7_inner_macOut <= _zz__16_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_518 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_6_inner_macOut;
  wire       [15:0]   _zz__zz__16_6_inner_macOut_1;
  wire       [15:0]   _zz__16_6_inner_macOut_1;
  wire       [15:0]   _zz__16_6_inner_macOut_2;
  reg        [7:0]    _16_6_inner_activation;
  reg        [7:0]    _16_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_6_inner_macOut;

  assign _zz__zz__16_6_inner_macOut = ($signed(io_mulInput) * $signed(_16_6_inner_activation));
  assign _zz__zz__16_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_6_inner_macOut)) ? 16'h007f : _zz__16_6_inner_macOut_2);
  assign _zz__16_6_inner_macOut_2 = (($signed(_zz__16_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_6_inner_activation;
    end else begin
      io_macOut = _16_6_inner_macOut;
    end
  end

  assign _zz__16_6_inner_macOut = ($signed(_zz__zz__16_6_inner_macOut) + $signed(_zz__zz__16_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_6_inner_activation <= 8'h00;
      _16_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_6_inner_activation <= io_addInput;
      end else begin
        _16_6_inner_macOut <= _zz__16_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_517 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_5_inner_macOut;
  wire       [15:0]   _zz__zz__16_5_inner_macOut_1;
  wire       [15:0]   _zz__16_5_inner_macOut_1;
  wire       [15:0]   _zz__16_5_inner_macOut_2;
  reg        [7:0]    _16_5_inner_activation;
  reg        [7:0]    _16_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_5_inner_macOut;

  assign _zz__zz__16_5_inner_macOut = ($signed(io_mulInput) * $signed(_16_5_inner_activation));
  assign _zz__zz__16_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_5_inner_macOut)) ? 16'h007f : _zz__16_5_inner_macOut_2);
  assign _zz__16_5_inner_macOut_2 = (($signed(_zz__16_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_5_inner_activation;
    end else begin
      io_macOut = _16_5_inner_macOut;
    end
  end

  assign _zz__16_5_inner_macOut = ($signed(_zz__zz__16_5_inner_macOut) + $signed(_zz__zz__16_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_5_inner_activation <= 8'h00;
      _16_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_5_inner_activation <= io_addInput;
      end else begin
        _16_5_inner_macOut <= _zz__16_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_516 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_4_inner_macOut;
  wire       [15:0]   _zz__zz__16_4_inner_macOut_1;
  wire       [15:0]   _zz__16_4_inner_macOut_1;
  wire       [15:0]   _zz__16_4_inner_macOut_2;
  reg        [7:0]    _16_4_inner_activation;
  reg        [7:0]    _16_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_4_inner_macOut;

  assign _zz__zz__16_4_inner_macOut = ($signed(io_mulInput) * $signed(_16_4_inner_activation));
  assign _zz__zz__16_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_4_inner_macOut)) ? 16'h007f : _zz__16_4_inner_macOut_2);
  assign _zz__16_4_inner_macOut_2 = (($signed(_zz__16_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_4_inner_activation;
    end else begin
      io_macOut = _16_4_inner_macOut;
    end
  end

  assign _zz__16_4_inner_macOut = ($signed(_zz__zz__16_4_inner_macOut) + $signed(_zz__zz__16_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_4_inner_activation <= 8'h00;
      _16_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_4_inner_activation <= io_addInput;
      end else begin
        _16_4_inner_macOut <= _zz__16_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_515 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_3_inner_macOut;
  wire       [15:0]   _zz__zz__16_3_inner_macOut_1;
  wire       [15:0]   _zz__16_3_inner_macOut_1;
  wire       [15:0]   _zz__16_3_inner_macOut_2;
  reg        [7:0]    _16_3_inner_activation;
  reg        [7:0]    _16_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_3_inner_macOut;

  assign _zz__zz__16_3_inner_macOut = ($signed(io_mulInput) * $signed(_16_3_inner_activation));
  assign _zz__zz__16_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_3_inner_macOut)) ? 16'h007f : _zz__16_3_inner_macOut_2);
  assign _zz__16_3_inner_macOut_2 = (($signed(_zz__16_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_3_inner_activation;
    end else begin
      io_macOut = _16_3_inner_macOut;
    end
  end

  assign _zz__16_3_inner_macOut = ($signed(_zz__zz__16_3_inner_macOut) + $signed(_zz__zz__16_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_3_inner_activation <= 8'h00;
      _16_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_3_inner_activation <= io_addInput;
      end else begin
        _16_3_inner_macOut <= _zz__16_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_514 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_2_inner_macOut;
  wire       [15:0]   _zz__zz__16_2_inner_macOut_1;
  wire       [15:0]   _zz__16_2_inner_macOut_1;
  wire       [15:0]   _zz__16_2_inner_macOut_2;
  reg        [7:0]    _16_2_inner_activation;
  reg        [7:0]    _16_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_2_inner_macOut;

  assign _zz__zz__16_2_inner_macOut = ($signed(io_mulInput) * $signed(_16_2_inner_activation));
  assign _zz__zz__16_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_2_inner_macOut)) ? 16'h007f : _zz__16_2_inner_macOut_2);
  assign _zz__16_2_inner_macOut_2 = (($signed(_zz__16_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_2_inner_activation;
    end else begin
      io_macOut = _16_2_inner_macOut;
    end
  end

  assign _zz__16_2_inner_macOut = ($signed(_zz__zz__16_2_inner_macOut) + $signed(_zz__zz__16_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_2_inner_activation <= 8'h00;
      _16_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_2_inner_activation <= io_addInput;
      end else begin
        _16_2_inner_macOut <= _zz__16_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_513 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_1_inner_macOut;
  wire       [15:0]   _zz__zz__16_1_inner_macOut_1;
  wire       [15:0]   _zz__16_1_inner_macOut_1;
  wire       [15:0]   _zz__16_1_inner_macOut_2;
  reg        [7:0]    _16_1_inner_activation;
  reg        [7:0]    _16_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_1_inner_macOut;

  assign _zz__zz__16_1_inner_macOut = ($signed(io_mulInput) * $signed(_16_1_inner_activation));
  assign _zz__zz__16_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_1_inner_macOut)) ? 16'h007f : _zz__16_1_inner_macOut_2);
  assign _zz__16_1_inner_macOut_2 = (($signed(_zz__16_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_1_inner_activation;
    end else begin
      io_macOut = _16_1_inner_macOut;
    end
  end

  assign _zz__16_1_inner_macOut = ($signed(_zz__zz__16_1_inner_macOut) + $signed(_zz__zz__16_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_1_inner_activation <= 8'h00;
      _16_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_1_inner_activation <= io_addInput;
      end else begin
        _16_1_inner_macOut <= _zz__16_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_512 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__16_0_inner_macOut;
  wire       [15:0]   _zz__zz__16_0_inner_macOut_1;
  wire       [15:0]   _zz__16_0_inner_macOut_1;
  wire       [15:0]   _zz__16_0_inner_macOut_2;
  reg        [7:0]    _16_0_inner_activation;
  reg        [7:0]    _16_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__16_0_inner_macOut;

  assign _zz__zz__16_0_inner_macOut = ($signed(io_mulInput) * $signed(_16_0_inner_activation));
  assign _zz__zz__16_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__16_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__16_0_inner_macOut)) ? 16'h007f : _zz__16_0_inner_macOut_2);
  assign _zz__16_0_inner_macOut_2 = (($signed(_zz__16_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__16_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _16_0_inner_activation;
    end else begin
      io_macOut = _16_0_inner_macOut;
    end
  end

  assign _zz__16_0_inner_macOut = ($signed(_zz__zz__16_0_inner_macOut) + $signed(_zz__zz__16_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _16_0_inner_activation <= 8'h00;
      _16_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _16_0_inner_activation <= io_addInput;
      end else begin
        _16_0_inner_macOut <= _zz__16_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_511 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_31_inner_macOut;
  wire       [15:0]   _zz__zz__15_31_inner_macOut_1;
  wire       [15:0]   _zz__15_31_inner_macOut_1;
  wire       [15:0]   _zz__15_31_inner_macOut_2;
  reg        [7:0]    _15_31_inner_activation;
  reg        [7:0]    _15_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_31_inner_macOut;

  assign _zz__zz__15_31_inner_macOut = ($signed(io_mulInput) * $signed(_15_31_inner_activation));
  assign _zz__zz__15_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_31_inner_macOut)) ? 16'h007f : _zz__15_31_inner_macOut_2);
  assign _zz__15_31_inner_macOut_2 = (($signed(_zz__15_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_31_inner_activation;
    end else begin
      io_macOut = _15_31_inner_macOut;
    end
  end

  assign _zz__15_31_inner_macOut = ($signed(_zz__zz__15_31_inner_macOut) + $signed(_zz__zz__15_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_31_inner_activation <= 8'h00;
      _15_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_31_inner_activation <= io_addInput;
      end else begin
        _15_31_inner_macOut <= _zz__15_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_510 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_30_inner_macOut;
  wire       [15:0]   _zz__zz__15_30_inner_macOut_1;
  wire       [15:0]   _zz__15_30_inner_macOut_1;
  wire       [15:0]   _zz__15_30_inner_macOut_2;
  reg        [7:0]    _15_30_inner_activation;
  reg        [7:0]    _15_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_30_inner_macOut;

  assign _zz__zz__15_30_inner_macOut = ($signed(io_mulInput) * $signed(_15_30_inner_activation));
  assign _zz__zz__15_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_30_inner_macOut)) ? 16'h007f : _zz__15_30_inner_macOut_2);
  assign _zz__15_30_inner_macOut_2 = (($signed(_zz__15_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_30_inner_activation;
    end else begin
      io_macOut = _15_30_inner_macOut;
    end
  end

  assign _zz__15_30_inner_macOut = ($signed(_zz__zz__15_30_inner_macOut) + $signed(_zz__zz__15_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_30_inner_activation <= 8'h00;
      _15_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_30_inner_activation <= io_addInput;
      end else begin
        _15_30_inner_macOut <= _zz__15_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_509 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_29_inner_macOut;
  wire       [15:0]   _zz__zz__15_29_inner_macOut_1;
  wire       [15:0]   _zz__15_29_inner_macOut_1;
  wire       [15:0]   _zz__15_29_inner_macOut_2;
  reg        [7:0]    _15_29_inner_activation;
  reg        [7:0]    _15_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_29_inner_macOut;

  assign _zz__zz__15_29_inner_macOut = ($signed(io_mulInput) * $signed(_15_29_inner_activation));
  assign _zz__zz__15_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_29_inner_macOut)) ? 16'h007f : _zz__15_29_inner_macOut_2);
  assign _zz__15_29_inner_macOut_2 = (($signed(_zz__15_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_29_inner_activation;
    end else begin
      io_macOut = _15_29_inner_macOut;
    end
  end

  assign _zz__15_29_inner_macOut = ($signed(_zz__zz__15_29_inner_macOut) + $signed(_zz__zz__15_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_29_inner_activation <= 8'h00;
      _15_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_29_inner_activation <= io_addInput;
      end else begin
        _15_29_inner_macOut <= _zz__15_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_508 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_28_inner_macOut;
  wire       [15:0]   _zz__zz__15_28_inner_macOut_1;
  wire       [15:0]   _zz__15_28_inner_macOut_1;
  wire       [15:0]   _zz__15_28_inner_macOut_2;
  reg        [7:0]    _15_28_inner_activation;
  reg        [7:0]    _15_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_28_inner_macOut;

  assign _zz__zz__15_28_inner_macOut = ($signed(io_mulInput) * $signed(_15_28_inner_activation));
  assign _zz__zz__15_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_28_inner_macOut)) ? 16'h007f : _zz__15_28_inner_macOut_2);
  assign _zz__15_28_inner_macOut_2 = (($signed(_zz__15_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_28_inner_activation;
    end else begin
      io_macOut = _15_28_inner_macOut;
    end
  end

  assign _zz__15_28_inner_macOut = ($signed(_zz__zz__15_28_inner_macOut) + $signed(_zz__zz__15_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_28_inner_activation <= 8'h00;
      _15_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_28_inner_activation <= io_addInput;
      end else begin
        _15_28_inner_macOut <= _zz__15_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_507 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_27_inner_macOut;
  wire       [15:0]   _zz__zz__15_27_inner_macOut_1;
  wire       [15:0]   _zz__15_27_inner_macOut_1;
  wire       [15:0]   _zz__15_27_inner_macOut_2;
  reg        [7:0]    _15_27_inner_activation;
  reg        [7:0]    _15_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_27_inner_macOut;

  assign _zz__zz__15_27_inner_macOut = ($signed(io_mulInput) * $signed(_15_27_inner_activation));
  assign _zz__zz__15_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_27_inner_macOut)) ? 16'h007f : _zz__15_27_inner_macOut_2);
  assign _zz__15_27_inner_macOut_2 = (($signed(_zz__15_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_27_inner_activation;
    end else begin
      io_macOut = _15_27_inner_macOut;
    end
  end

  assign _zz__15_27_inner_macOut = ($signed(_zz__zz__15_27_inner_macOut) + $signed(_zz__zz__15_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_27_inner_activation <= 8'h00;
      _15_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_27_inner_activation <= io_addInput;
      end else begin
        _15_27_inner_macOut <= _zz__15_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_506 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_26_inner_macOut;
  wire       [15:0]   _zz__zz__15_26_inner_macOut_1;
  wire       [15:0]   _zz__15_26_inner_macOut_1;
  wire       [15:0]   _zz__15_26_inner_macOut_2;
  reg        [7:0]    _15_26_inner_activation;
  reg        [7:0]    _15_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_26_inner_macOut;

  assign _zz__zz__15_26_inner_macOut = ($signed(io_mulInput) * $signed(_15_26_inner_activation));
  assign _zz__zz__15_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_26_inner_macOut)) ? 16'h007f : _zz__15_26_inner_macOut_2);
  assign _zz__15_26_inner_macOut_2 = (($signed(_zz__15_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_26_inner_activation;
    end else begin
      io_macOut = _15_26_inner_macOut;
    end
  end

  assign _zz__15_26_inner_macOut = ($signed(_zz__zz__15_26_inner_macOut) + $signed(_zz__zz__15_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_26_inner_activation <= 8'h00;
      _15_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_26_inner_activation <= io_addInput;
      end else begin
        _15_26_inner_macOut <= _zz__15_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_505 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_25_inner_macOut;
  wire       [15:0]   _zz__zz__15_25_inner_macOut_1;
  wire       [15:0]   _zz__15_25_inner_macOut_1;
  wire       [15:0]   _zz__15_25_inner_macOut_2;
  reg        [7:0]    _15_25_inner_activation;
  reg        [7:0]    _15_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_25_inner_macOut;

  assign _zz__zz__15_25_inner_macOut = ($signed(io_mulInput) * $signed(_15_25_inner_activation));
  assign _zz__zz__15_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_25_inner_macOut)) ? 16'h007f : _zz__15_25_inner_macOut_2);
  assign _zz__15_25_inner_macOut_2 = (($signed(_zz__15_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_25_inner_activation;
    end else begin
      io_macOut = _15_25_inner_macOut;
    end
  end

  assign _zz__15_25_inner_macOut = ($signed(_zz__zz__15_25_inner_macOut) + $signed(_zz__zz__15_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_25_inner_activation <= 8'h00;
      _15_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_25_inner_activation <= io_addInput;
      end else begin
        _15_25_inner_macOut <= _zz__15_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_504 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_24_inner_macOut;
  wire       [15:0]   _zz__zz__15_24_inner_macOut_1;
  wire       [15:0]   _zz__15_24_inner_macOut_1;
  wire       [15:0]   _zz__15_24_inner_macOut_2;
  reg        [7:0]    _15_24_inner_activation;
  reg        [7:0]    _15_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_24_inner_macOut;

  assign _zz__zz__15_24_inner_macOut = ($signed(io_mulInput) * $signed(_15_24_inner_activation));
  assign _zz__zz__15_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_24_inner_macOut)) ? 16'h007f : _zz__15_24_inner_macOut_2);
  assign _zz__15_24_inner_macOut_2 = (($signed(_zz__15_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_24_inner_activation;
    end else begin
      io_macOut = _15_24_inner_macOut;
    end
  end

  assign _zz__15_24_inner_macOut = ($signed(_zz__zz__15_24_inner_macOut) + $signed(_zz__zz__15_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_24_inner_activation <= 8'h00;
      _15_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_24_inner_activation <= io_addInput;
      end else begin
        _15_24_inner_macOut <= _zz__15_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_503 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_23_inner_macOut;
  wire       [15:0]   _zz__zz__15_23_inner_macOut_1;
  wire       [15:0]   _zz__15_23_inner_macOut_1;
  wire       [15:0]   _zz__15_23_inner_macOut_2;
  reg        [7:0]    _15_23_inner_activation;
  reg        [7:0]    _15_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_23_inner_macOut;

  assign _zz__zz__15_23_inner_macOut = ($signed(io_mulInput) * $signed(_15_23_inner_activation));
  assign _zz__zz__15_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_23_inner_macOut)) ? 16'h007f : _zz__15_23_inner_macOut_2);
  assign _zz__15_23_inner_macOut_2 = (($signed(_zz__15_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_23_inner_activation;
    end else begin
      io_macOut = _15_23_inner_macOut;
    end
  end

  assign _zz__15_23_inner_macOut = ($signed(_zz__zz__15_23_inner_macOut) + $signed(_zz__zz__15_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_23_inner_activation <= 8'h00;
      _15_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_23_inner_activation <= io_addInput;
      end else begin
        _15_23_inner_macOut <= _zz__15_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_502 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_22_inner_macOut;
  wire       [15:0]   _zz__zz__15_22_inner_macOut_1;
  wire       [15:0]   _zz__15_22_inner_macOut_1;
  wire       [15:0]   _zz__15_22_inner_macOut_2;
  reg        [7:0]    _15_22_inner_activation;
  reg        [7:0]    _15_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_22_inner_macOut;

  assign _zz__zz__15_22_inner_macOut = ($signed(io_mulInput) * $signed(_15_22_inner_activation));
  assign _zz__zz__15_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_22_inner_macOut)) ? 16'h007f : _zz__15_22_inner_macOut_2);
  assign _zz__15_22_inner_macOut_2 = (($signed(_zz__15_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_22_inner_activation;
    end else begin
      io_macOut = _15_22_inner_macOut;
    end
  end

  assign _zz__15_22_inner_macOut = ($signed(_zz__zz__15_22_inner_macOut) + $signed(_zz__zz__15_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_22_inner_activation <= 8'h00;
      _15_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_22_inner_activation <= io_addInput;
      end else begin
        _15_22_inner_macOut <= _zz__15_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_501 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_21_inner_macOut;
  wire       [15:0]   _zz__zz__15_21_inner_macOut_1;
  wire       [15:0]   _zz__15_21_inner_macOut_1;
  wire       [15:0]   _zz__15_21_inner_macOut_2;
  reg        [7:0]    _15_21_inner_activation;
  reg        [7:0]    _15_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_21_inner_macOut;

  assign _zz__zz__15_21_inner_macOut = ($signed(io_mulInput) * $signed(_15_21_inner_activation));
  assign _zz__zz__15_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_21_inner_macOut)) ? 16'h007f : _zz__15_21_inner_macOut_2);
  assign _zz__15_21_inner_macOut_2 = (($signed(_zz__15_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_21_inner_activation;
    end else begin
      io_macOut = _15_21_inner_macOut;
    end
  end

  assign _zz__15_21_inner_macOut = ($signed(_zz__zz__15_21_inner_macOut) + $signed(_zz__zz__15_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_21_inner_activation <= 8'h00;
      _15_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_21_inner_activation <= io_addInput;
      end else begin
        _15_21_inner_macOut <= _zz__15_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_500 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_20_inner_macOut;
  wire       [15:0]   _zz__zz__15_20_inner_macOut_1;
  wire       [15:0]   _zz__15_20_inner_macOut_1;
  wire       [15:0]   _zz__15_20_inner_macOut_2;
  reg        [7:0]    _15_20_inner_activation;
  reg        [7:0]    _15_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_20_inner_macOut;

  assign _zz__zz__15_20_inner_macOut = ($signed(io_mulInput) * $signed(_15_20_inner_activation));
  assign _zz__zz__15_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_20_inner_macOut)) ? 16'h007f : _zz__15_20_inner_macOut_2);
  assign _zz__15_20_inner_macOut_2 = (($signed(_zz__15_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_20_inner_activation;
    end else begin
      io_macOut = _15_20_inner_macOut;
    end
  end

  assign _zz__15_20_inner_macOut = ($signed(_zz__zz__15_20_inner_macOut) + $signed(_zz__zz__15_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_20_inner_activation <= 8'h00;
      _15_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_20_inner_activation <= io_addInput;
      end else begin
        _15_20_inner_macOut <= _zz__15_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_499 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_19_inner_macOut;
  wire       [15:0]   _zz__zz__15_19_inner_macOut_1;
  wire       [15:0]   _zz__15_19_inner_macOut_1;
  wire       [15:0]   _zz__15_19_inner_macOut_2;
  reg        [7:0]    _15_19_inner_activation;
  reg        [7:0]    _15_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_19_inner_macOut;

  assign _zz__zz__15_19_inner_macOut = ($signed(io_mulInput) * $signed(_15_19_inner_activation));
  assign _zz__zz__15_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_19_inner_macOut)) ? 16'h007f : _zz__15_19_inner_macOut_2);
  assign _zz__15_19_inner_macOut_2 = (($signed(_zz__15_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_19_inner_activation;
    end else begin
      io_macOut = _15_19_inner_macOut;
    end
  end

  assign _zz__15_19_inner_macOut = ($signed(_zz__zz__15_19_inner_macOut) + $signed(_zz__zz__15_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_19_inner_activation <= 8'h00;
      _15_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_19_inner_activation <= io_addInput;
      end else begin
        _15_19_inner_macOut <= _zz__15_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_498 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_18_inner_macOut;
  wire       [15:0]   _zz__zz__15_18_inner_macOut_1;
  wire       [15:0]   _zz__15_18_inner_macOut_1;
  wire       [15:0]   _zz__15_18_inner_macOut_2;
  reg        [7:0]    _15_18_inner_activation;
  reg        [7:0]    _15_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_18_inner_macOut;

  assign _zz__zz__15_18_inner_macOut = ($signed(io_mulInput) * $signed(_15_18_inner_activation));
  assign _zz__zz__15_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_18_inner_macOut)) ? 16'h007f : _zz__15_18_inner_macOut_2);
  assign _zz__15_18_inner_macOut_2 = (($signed(_zz__15_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_18_inner_activation;
    end else begin
      io_macOut = _15_18_inner_macOut;
    end
  end

  assign _zz__15_18_inner_macOut = ($signed(_zz__zz__15_18_inner_macOut) + $signed(_zz__zz__15_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_18_inner_activation <= 8'h00;
      _15_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_18_inner_activation <= io_addInput;
      end else begin
        _15_18_inner_macOut <= _zz__15_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_497 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_17_inner_macOut;
  wire       [15:0]   _zz__zz__15_17_inner_macOut_1;
  wire       [15:0]   _zz__15_17_inner_macOut_1;
  wire       [15:0]   _zz__15_17_inner_macOut_2;
  reg        [7:0]    _15_17_inner_activation;
  reg        [7:0]    _15_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_17_inner_macOut;

  assign _zz__zz__15_17_inner_macOut = ($signed(io_mulInput) * $signed(_15_17_inner_activation));
  assign _zz__zz__15_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_17_inner_macOut)) ? 16'h007f : _zz__15_17_inner_macOut_2);
  assign _zz__15_17_inner_macOut_2 = (($signed(_zz__15_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_17_inner_activation;
    end else begin
      io_macOut = _15_17_inner_macOut;
    end
  end

  assign _zz__15_17_inner_macOut = ($signed(_zz__zz__15_17_inner_macOut) + $signed(_zz__zz__15_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_17_inner_activation <= 8'h00;
      _15_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_17_inner_activation <= io_addInput;
      end else begin
        _15_17_inner_macOut <= _zz__15_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_496 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_16_inner_macOut;
  wire       [15:0]   _zz__zz__15_16_inner_macOut_1;
  wire       [15:0]   _zz__15_16_inner_macOut_1;
  wire       [15:0]   _zz__15_16_inner_macOut_2;
  reg        [7:0]    _15_16_inner_activation;
  reg        [7:0]    _15_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_16_inner_macOut;

  assign _zz__zz__15_16_inner_macOut = ($signed(io_mulInput) * $signed(_15_16_inner_activation));
  assign _zz__zz__15_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_16_inner_macOut)) ? 16'h007f : _zz__15_16_inner_macOut_2);
  assign _zz__15_16_inner_macOut_2 = (($signed(_zz__15_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_16_inner_activation;
    end else begin
      io_macOut = _15_16_inner_macOut;
    end
  end

  assign _zz__15_16_inner_macOut = ($signed(_zz__zz__15_16_inner_macOut) + $signed(_zz__zz__15_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_16_inner_activation <= 8'h00;
      _15_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_16_inner_activation <= io_addInput;
      end else begin
        _15_16_inner_macOut <= _zz__15_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_495 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_15_inner_macOut;
  wire       [15:0]   _zz__zz__15_15_inner_macOut_1;
  wire       [15:0]   _zz__15_15_inner_macOut_1;
  wire       [15:0]   _zz__15_15_inner_macOut_2;
  reg        [7:0]    _15_15_inner_activation;
  reg        [7:0]    _15_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_15_inner_macOut;

  assign _zz__zz__15_15_inner_macOut = ($signed(io_mulInput) * $signed(_15_15_inner_activation));
  assign _zz__zz__15_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_15_inner_macOut)) ? 16'h007f : _zz__15_15_inner_macOut_2);
  assign _zz__15_15_inner_macOut_2 = (($signed(_zz__15_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_15_inner_activation;
    end else begin
      io_macOut = _15_15_inner_macOut;
    end
  end

  assign _zz__15_15_inner_macOut = ($signed(_zz__zz__15_15_inner_macOut) + $signed(_zz__zz__15_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_15_inner_activation <= 8'h00;
      _15_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_15_inner_activation <= io_addInput;
      end else begin
        _15_15_inner_macOut <= _zz__15_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_494 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_14_inner_macOut;
  wire       [15:0]   _zz__zz__15_14_inner_macOut_1;
  wire       [15:0]   _zz__15_14_inner_macOut_1;
  wire       [15:0]   _zz__15_14_inner_macOut_2;
  reg        [7:0]    _15_14_inner_activation;
  reg        [7:0]    _15_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_14_inner_macOut;

  assign _zz__zz__15_14_inner_macOut = ($signed(io_mulInput) * $signed(_15_14_inner_activation));
  assign _zz__zz__15_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_14_inner_macOut)) ? 16'h007f : _zz__15_14_inner_macOut_2);
  assign _zz__15_14_inner_macOut_2 = (($signed(_zz__15_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_14_inner_activation;
    end else begin
      io_macOut = _15_14_inner_macOut;
    end
  end

  assign _zz__15_14_inner_macOut = ($signed(_zz__zz__15_14_inner_macOut) + $signed(_zz__zz__15_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_14_inner_activation <= 8'h00;
      _15_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_14_inner_activation <= io_addInput;
      end else begin
        _15_14_inner_macOut <= _zz__15_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_493 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_13_inner_macOut;
  wire       [15:0]   _zz__zz__15_13_inner_macOut_1;
  wire       [15:0]   _zz__15_13_inner_macOut_1;
  wire       [15:0]   _zz__15_13_inner_macOut_2;
  reg        [7:0]    _15_13_inner_activation;
  reg        [7:0]    _15_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_13_inner_macOut;

  assign _zz__zz__15_13_inner_macOut = ($signed(io_mulInput) * $signed(_15_13_inner_activation));
  assign _zz__zz__15_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_13_inner_macOut)) ? 16'h007f : _zz__15_13_inner_macOut_2);
  assign _zz__15_13_inner_macOut_2 = (($signed(_zz__15_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_13_inner_activation;
    end else begin
      io_macOut = _15_13_inner_macOut;
    end
  end

  assign _zz__15_13_inner_macOut = ($signed(_zz__zz__15_13_inner_macOut) + $signed(_zz__zz__15_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_13_inner_activation <= 8'h00;
      _15_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_13_inner_activation <= io_addInput;
      end else begin
        _15_13_inner_macOut <= _zz__15_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_492 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_12_inner_macOut;
  wire       [15:0]   _zz__zz__15_12_inner_macOut_1;
  wire       [15:0]   _zz__15_12_inner_macOut_1;
  wire       [15:0]   _zz__15_12_inner_macOut_2;
  reg        [7:0]    _15_12_inner_activation;
  reg        [7:0]    _15_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_12_inner_macOut;

  assign _zz__zz__15_12_inner_macOut = ($signed(io_mulInput) * $signed(_15_12_inner_activation));
  assign _zz__zz__15_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_12_inner_macOut)) ? 16'h007f : _zz__15_12_inner_macOut_2);
  assign _zz__15_12_inner_macOut_2 = (($signed(_zz__15_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_12_inner_activation;
    end else begin
      io_macOut = _15_12_inner_macOut;
    end
  end

  assign _zz__15_12_inner_macOut = ($signed(_zz__zz__15_12_inner_macOut) + $signed(_zz__zz__15_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_12_inner_activation <= 8'h00;
      _15_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_12_inner_activation <= io_addInput;
      end else begin
        _15_12_inner_macOut <= _zz__15_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_491 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_11_inner_macOut;
  wire       [15:0]   _zz__zz__15_11_inner_macOut_1;
  wire       [15:0]   _zz__15_11_inner_macOut_1;
  wire       [15:0]   _zz__15_11_inner_macOut_2;
  reg        [7:0]    _15_11_inner_activation;
  reg        [7:0]    _15_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_11_inner_macOut;

  assign _zz__zz__15_11_inner_macOut = ($signed(io_mulInput) * $signed(_15_11_inner_activation));
  assign _zz__zz__15_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_11_inner_macOut)) ? 16'h007f : _zz__15_11_inner_macOut_2);
  assign _zz__15_11_inner_macOut_2 = (($signed(_zz__15_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_11_inner_activation;
    end else begin
      io_macOut = _15_11_inner_macOut;
    end
  end

  assign _zz__15_11_inner_macOut = ($signed(_zz__zz__15_11_inner_macOut) + $signed(_zz__zz__15_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_11_inner_activation <= 8'h00;
      _15_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_11_inner_activation <= io_addInput;
      end else begin
        _15_11_inner_macOut <= _zz__15_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_490 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_10_inner_macOut;
  wire       [15:0]   _zz__zz__15_10_inner_macOut_1;
  wire       [15:0]   _zz__15_10_inner_macOut_1;
  wire       [15:0]   _zz__15_10_inner_macOut_2;
  reg        [7:0]    _15_10_inner_activation;
  reg        [7:0]    _15_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_10_inner_macOut;

  assign _zz__zz__15_10_inner_macOut = ($signed(io_mulInput) * $signed(_15_10_inner_activation));
  assign _zz__zz__15_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_10_inner_macOut)) ? 16'h007f : _zz__15_10_inner_macOut_2);
  assign _zz__15_10_inner_macOut_2 = (($signed(_zz__15_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_10_inner_activation;
    end else begin
      io_macOut = _15_10_inner_macOut;
    end
  end

  assign _zz__15_10_inner_macOut = ($signed(_zz__zz__15_10_inner_macOut) + $signed(_zz__zz__15_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_10_inner_activation <= 8'h00;
      _15_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_10_inner_activation <= io_addInput;
      end else begin
        _15_10_inner_macOut <= _zz__15_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_489 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_9_inner_macOut;
  wire       [15:0]   _zz__zz__15_9_inner_macOut_1;
  wire       [15:0]   _zz__15_9_inner_macOut_1;
  wire       [15:0]   _zz__15_9_inner_macOut_2;
  reg        [7:0]    _15_9_inner_activation;
  reg        [7:0]    _15_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_9_inner_macOut;

  assign _zz__zz__15_9_inner_macOut = ($signed(io_mulInput) * $signed(_15_9_inner_activation));
  assign _zz__zz__15_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_9_inner_macOut)) ? 16'h007f : _zz__15_9_inner_macOut_2);
  assign _zz__15_9_inner_macOut_2 = (($signed(_zz__15_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_9_inner_activation;
    end else begin
      io_macOut = _15_9_inner_macOut;
    end
  end

  assign _zz__15_9_inner_macOut = ($signed(_zz__zz__15_9_inner_macOut) + $signed(_zz__zz__15_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_9_inner_activation <= 8'h00;
      _15_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_9_inner_activation <= io_addInput;
      end else begin
        _15_9_inner_macOut <= _zz__15_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_488 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_8_inner_macOut;
  wire       [15:0]   _zz__zz__15_8_inner_macOut_1;
  wire       [15:0]   _zz__15_8_inner_macOut_1;
  wire       [15:0]   _zz__15_8_inner_macOut_2;
  reg        [7:0]    _15_8_inner_activation;
  reg        [7:0]    _15_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_8_inner_macOut;

  assign _zz__zz__15_8_inner_macOut = ($signed(io_mulInput) * $signed(_15_8_inner_activation));
  assign _zz__zz__15_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_8_inner_macOut)) ? 16'h007f : _zz__15_8_inner_macOut_2);
  assign _zz__15_8_inner_macOut_2 = (($signed(_zz__15_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_8_inner_activation;
    end else begin
      io_macOut = _15_8_inner_macOut;
    end
  end

  assign _zz__15_8_inner_macOut = ($signed(_zz__zz__15_8_inner_macOut) + $signed(_zz__zz__15_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_8_inner_activation <= 8'h00;
      _15_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_8_inner_activation <= io_addInput;
      end else begin
        _15_8_inner_macOut <= _zz__15_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_487 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_7_inner_macOut;
  wire       [15:0]   _zz__zz__15_7_inner_macOut_1;
  wire       [15:0]   _zz__15_7_inner_macOut_1;
  wire       [15:0]   _zz__15_7_inner_macOut_2;
  reg        [7:0]    _15_7_inner_activation;
  reg        [7:0]    _15_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_7_inner_macOut;

  assign _zz__zz__15_7_inner_macOut = ($signed(io_mulInput) * $signed(_15_7_inner_activation));
  assign _zz__zz__15_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_7_inner_macOut)) ? 16'h007f : _zz__15_7_inner_macOut_2);
  assign _zz__15_7_inner_macOut_2 = (($signed(_zz__15_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_7_inner_activation;
    end else begin
      io_macOut = _15_7_inner_macOut;
    end
  end

  assign _zz__15_7_inner_macOut = ($signed(_zz__zz__15_7_inner_macOut) + $signed(_zz__zz__15_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_7_inner_activation <= 8'h00;
      _15_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_7_inner_activation <= io_addInput;
      end else begin
        _15_7_inner_macOut <= _zz__15_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_486 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_6_inner_macOut;
  wire       [15:0]   _zz__zz__15_6_inner_macOut_1;
  wire       [15:0]   _zz__15_6_inner_macOut_1;
  wire       [15:0]   _zz__15_6_inner_macOut_2;
  reg        [7:0]    _15_6_inner_activation;
  reg        [7:0]    _15_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_6_inner_macOut;

  assign _zz__zz__15_6_inner_macOut = ($signed(io_mulInput) * $signed(_15_6_inner_activation));
  assign _zz__zz__15_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_6_inner_macOut)) ? 16'h007f : _zz__15_6_inner_macOut_2);
  assign _zz__15_6_inner_macOut_2 = (($signed(_zz__15_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_6_inner_activation;
    end else begin
      io_macOut = _15_6_inner_macOut;
    end
  end

  assign _zz__15_6_inner_macOut = ($signed(_zz__zz__15_6_inner_macOut) + $signed(_zz__zz__15_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_6_inner_activation <= 8'h00;
      _15_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_6_inner_activation <= io_addInput;
      end else begin
        _15_6_inner_macOut <= _zz__15_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_485 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_5_inner_macOut;
  wire       [15:0]   _zz__zz__15_5_inner_macOut_1;
  wire       [15:0]   _zz__15_5_inner_macOut_1;
  wire       [15:0]   _zz__15_5_inner_macOut_2;
  reg        [7:0]    _15_5_inner_activation;
  reg        [7:0]    _15_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_5_inner_macOut;

  assign _zz__zz__15_5_inner_macOut = ($signed(io_mulInput) * $signed(_15_5_inner_activation));
  assign _zz__zz__15_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_5_inner_macOut)) ? 16'h007f : _zz__15_5_inner_macOut_2);
  assign _zz__15_5_inner_macOut_2 = (($signed(_zz__15_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_5_inner_activation;
    end else begin
      io_macOut = _15_5_inner_macOut;
    end
  end

  assign _zz__15_5_inner_macOut = ($signed(_zz__zz__15_5_inner_macOut) + $signed(_zz__zz__15_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_5_inner_activation <= 8'h00;
      _15_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_5_inner_activation <= io_addInput;
      end else begin
        _15_5_inner_macOut <= _zz__15_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_484 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_4_inner_macOut;
  wire       [15:0]   _zz__zz__15_4_inner_macOut_1;
  wire       [15:0]   _zz__15_4_inner_macOut_1;
  wire       [15:0]   _zz__15_4_inner_macOut_2;
  reg        [7:0]    _15_4_inner_activation;
  reg        [7:0]    _15_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_4_inner_macOut;

  assign _zz__zz__15_4_inner_macOut = ($signed(io_mulInput) * $signed(_15_4_inner_activation));
  assign _zz__zz__15_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_4_inner_macOut)) ? 16'h007f : _zz__15_4_inner_macOut_2);
  assign _zz__15_4_inner_macOut_2 = (($signed(_zz__15_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_4_inner_activation;
    end else begin
      io_macOut = _15_4_inner_macOut;
    end
  end

  assign _zz__15_4_inner_macOut = ($signed(_zz__zz__15_4_inner_macOut) + $signed(_zz__zz__15_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_4_inner_activation <= 8'h00;
      _15_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_4_inner_activation <= io_addInput;
      end else begin
        _15_4_inner_macOut <= _zz__15_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_483 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_3_inner_macOut;
  wire       [15:0]   _zz__zz__15_3_inner_macOut_1;
  wire       [15:0]   _zz__15_3_inner_macOut_1;
  wire       [15:0]   _zz__15_3_inner_macOut_2;
  reg        [7:0]    _15_3_inner_activation;
  reg        [7:0]    _15_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_3_inner_macOut;

  assign _zz__zz__15_3_inner_macOut = ($signed(io_mulInput) * $signed(_15_3_inner_activation));
  assign _zz__zz__15_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_3_inner_macOut)) ? 16'h007f : _zz__15_3_inner_macOut_2);
  assign _zz__15_3_inner_macOut_2 = (($signed(_zz__15_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_3_inner_activation;
    end else begin
      io_macOut = _15_3_inner_macOut;
    end
  end

  assign _zz__15_3_inner_macOut = ($signed(_zz__zz__15_3_inner_macOut) + $signed(_zz__zz__15_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_3_inner_activation <= 8'h00;
      _15_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_3_inner_activation <= io_addInput;
      end else begin
        _15_3_inner_macOut <= _zz__15_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_482 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_2_inner_macOut;
  wire       [15:0]   _zz__zz__15_2_inner_macOut_1;
  wire       [15:0]   _zz__15_2_inner_macOut_1;
  wire       [15:0]   _zz__15_2_inner_macOut_2;
  reg        [7:0]    _15_2_inner_activation;
  reg        [7:0]    _15_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_2_inner_macOut;

  assign _zz__zz__15_2_inner_macOut = ($signed(io_mulInput) * $signed(_15_2_inner_activation));
  assign _zz__zz__15_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_2_inner_macOut)) ? 16'h007f : _zz__15_2_inner_macOut_2);
  assign _zz__15_2_inner_macOut_2 = (($signed(_zz__15_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_2_inner_activation;
    end else begin
      io_macOut = _15_2_inner_macOut;
    end
  end

  assign _zz__15_2_inner_macOut = ($signed(_zz__zz__15_2_inner_macOut) + $signed(_zz__zz__15_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_2_inner_activation <= 8'h00;
      _15_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_2_inner_activation <= io_addInput;
      end else begin
        _15_2_inner_macOut <= _zz__15_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_481 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_1_inner_macOut;
  wire       [15:0]   _zz__zz__15_1_inner_macOut_1;
  wire       [15:0]   _zz__15_1_inner_macOut_1;
  wire       [15:0]   _zz__15_1_inner_macOut_2;
  reg        [7:0]    _15_1_inner_activation;
  reg        [7:0]    _15_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_1_inner_macOut;

  assign _zz__zz__15_1_inner_macOut = ($signed(io_mulInput) * $signed(_15_1_inner_activation));
  assign _zz__zz__15_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_1_inner_macOut)) ? 16'h007f : _zz__15_1_inner_macOut_2);
  assign _zz__15_1_inner_macOut_2 = (($signed(_zz__15_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_1_inner_activation;
    end else begin
      io_macOut = _15_1_inner_macOut;
    end
  end

  assign _zz__15_1_inner_macOut = ($signed(_zz__zz__15_1_inner_macOut) + $signed(_zz__zz__15_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_1_inner_activation <= 8'h00;
      _15_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_1_inner_activation <= io_addInput;
      end else begin
        _15_1_inner_macOut <= _zz__15_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_480 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__15_0_inner_macOut;
  wire       [15:0]   _zz__zz__15_0_inner_macOut_1;
  wire       [15:0]   _zz__15_0_inner_macOut_1;
  wire       [15:0]   _zz__15_0_inner_macOut_2;
  reg        [7:0]    _15_0_inner_activation;
  reg        [7:0]    _15_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__15_0_inner_macOut;

  assign _zz__zz__15_0_inner_macOut = ($signed(io_mulInput) * $signed(_15_0_inner_activation));
  assign _zz__zz__15_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__15_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__15_0_inner_macOut)) ? 16'h007f : _zz__15_0_inner_macOut_2);
  assign _zz__15_0_inner_macOut_2 = (($signed(_zz__15_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__15_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _15_0_inner_activation;
    end else begin
      io_macOut = _15_0_inner_macOut;
    end
  end

  assign _zz__15_0_inner_macOut = ($signed(_zz__zz__15_0_inner_macOut) + $signed(_zz__zz__15_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _15_0_inner_activation <= 8'h00;
      _15_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _15_0_inner_activation <= io_addInput;
      end else begin
        _15_0_inner_macOut <= _zz__15_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_479 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_31_inner_macOut;
  wire       [15:0]   _zz__zz__14_31_inner_macOut_1;
  wire       [15:0]   _zz__14_31_inner_macOut_1;
  wire       [15:0]   _zz__14_31_inner_macOut_2;
  reg        [7:0]    _14_31_inner_activation;
  reg        [7:0]    _14_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_31_inner_macOut;

  assign _zz__zz__14_31_inner_macOut = ($signed(io_mulInput) * $signed(_14_31_inner_activation));
  assign _zz__zz__14_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_31_inner_macOut)) ? 16'h007f : _zz__14_31_inner_macOut_2);
  assign _zz__14_31_inner_macOut_2 = (($signed(_zz__14_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_31_inner_activation;
    end else begin
      io_macOut = _14_31_inner_macOut;
    end
  end

  assign _zz__14_31_inner_macOut = ($signed(_zz__zz__14_31_inner_macOut) + $signed(_zz__zz__14_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_31_inner_activation <= 8'h00;
      _14_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_31_inner_activation <= io_addInput;
      end else begin
        _14_31_inner_macOut <= _zz__14_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_478 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_30_inner_macOut;
  wire       [15:0]   _zz__zz__14_30_inner_macOut_1;
  wire       [15:0]   _zz__14_30_inner_macOut_1;
  wire       [15:0]   _zz__14_30_inner_macOut_2;
  reg        [7:0]    _14_30_inner_activation;
  reg        [7:0]    _14_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_30_inner_macOut;

  assign _zz__zz__14_30_inner_macOut = ($signed(io_mulInput) * $signed(_14_30_inner_activation));
  assign _zz__zz__14_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_30_inner_macOut)) ? 16'h007f : _zz__14_30_inner_macOut_2);
  assign _zz__14_30_inner_macOut_2 = (($signed(_zz__14_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_30_inner_activation;
    end else begin
      io_macOut = _14_30_inner_macOut;
    end
  end

  assign _zz__14_30_inner_macOut = ($signed(_zz__zz__14_30_inner_macOut) + $signed(_zz__zz__14_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_30_inner_activation <= 8'h00;
      _14_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_30_inner_activation <= io_addInput;
      end else begin
        _14_30_inner_macOut <= _zz__14_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_477 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_29_inner_macOut;
  wire       [15:0]   _zz__zz__14_29_inner_macOut_1;
  wire       [15:0]   _zz__14_29_inner_macOut_1;
  wire       [15:0]   _zz__14_29_inner_macOut_2;
  reg        [7:0]    _14_29_inner_activation;
  reg        [7:0]    _14_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_29_inner_macOut;

  assign _zz__zz__14_29_inner_macOut = ($signed(io_mulInput) * $signed(_14_29_inner_activation));
  assign _zz__zz__14_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_29_inner_macOut)) ? 16'h007f : _zz__14_29_inner_macOut_2);
  assign _zz__14_29_inner_macOut_2 = (($signed(_zz__14_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_29_inner_activation;
    end else begin
      io_macOut = _14_29_inner_macOut;
    end
  end

  assign _zz__14_29_inner_macOut = ($signed(_zz__zz__14_29_inner_macOut) + $signed(_zz__zz__14_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_29_inner_activation <= 8'h00;
      _14_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_29_inner_activation <= io_addInput;
      end else begin
        _14_29_inner_macOut <= _zz__14_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_476 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_28_inner_macOut;
  wire       [15:0]   _zz__zz__14_28_inner_macOut_1;
  wire       [15:0]   _zz__14_28_inner_macOut_1;
  wire       [15:0]   _zz__14_28_inner_macOut_2;
  reg        [7:0]    _14_28_inner_activation;
  reg        [7:0]    _14_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_28_inner_macOut;

  assign _zz__zz__14_28_inner_macOut = ($signed(io_mulInput) * $signed(_14_28_inner_activation));
  assign _zz__zz__14_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_28_inner_macOut)) ? 16'h007f : _zz__14_28_inner_macOut_2);
  assign _zz__14_28_inner_macOut_2 = (($signed(_zz__14_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_28_inner_activation;
    end else begin
      io_macOut = _14_28_inner_macOut;
    end
  end

  assign _zz__14_28_inner_macOut = ($signed(_zz__zz__14_28_inner_macOut) + $signed(_zz__zz__14_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_28_inner_activation <= 8'h00;
      _14_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_28_inner_activation <= io_addInput;
      end else begin
        _14_28_inner_macOut <= _zz__14_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_475 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_27_inner_macOut;
  wire       [15:0]   _zz__zz__14_27_inner_macOut_1;
  wire       [15:0]   _zz__14_27_inner_macOut_1;
  wire       [15:0]   _zz__14_27_inner_macOut_2;
  reg        [7:0]    _14_27_inner_activation;
  reg        [7:0]    _14_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_27_inner_macOut;

  assign _zz__zz__14_27_inner_macOut = ($signed(io_mulInput) * $signed(_14_27_inner_activation));
  assign _zz__zz__14_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_27_inner_macOut)) ? 16'h007f : _zz__14_27_inner_macOut_2);
  assign _zz__14_27_inner_macOut_2 = (($signed(_zz__14_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_27_inner_activation;
    end else begin
      io_macOut = _14_27_inner_macOut;
    end
  end

  assign _zz__14_27_inner_macOut = ($signed(_zz__zz__14_27_inner_macOut) + $signed(_zz__zz__14_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_27_inner_activation <= 8'h00;
      _14_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_27_inner_activation <= io_addInput;
      end else begin
        _14_27_inner_macOut <= _zz__14_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_474 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_26_inner_macOut;
  wire       [15:0]   _zz__zz__14_26_inner_macOut_1;
  wire       [15:0]   _zz__14_26_inner_macOut_1;
  wire       [15:0]   _zz__14_26_inner_macOut_2;
  reg        [7:0]    _14_26_inner_activation;
  reg        [7:0]    _14_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_26_inner_macOut;

  assign _zz__zz__14_26_inner_macOut = ($signed(io_mulInput) * $signed(_14_26_inner_activation));
  assign _zz__zz__14_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_26_inner_macOut)) ? 16'h007f : _zz__14_26_inner_macOut_2);
  assign _zz__14_26_inner_macOut_2 = (($signed(_zz__14_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_26_inner_activation;
    end else begin
      io_macOut = _14_26_inner_macOut;
    end
  end

  assign _zz__14_26_inner_macOut = ($signed(_zz__zz__14_26_inner_macOut) + $signed(_zz__zz__14_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_26_inner_activation <= 8'h00;
      _14_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_26_inner_activation <= io_addInput;
      end else begin
        _14_26_inner_macOut <= _zz__14_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_473 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_25_inner_macOut;
  wire       [15:0]   _zz__zz__14_25_inner_macOut_1;
  wire       [15:0]   _zz__14_25_inner_macOut_1;
  wire       [15:0]   _zz__14_25_inner_macOut_2;
  reg        [7:0]    _14_25_inner_activation;
  reg        [7:0]    _14_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_25_inner_macOut;

  assign _zz__zz__14_25_inner_macOut = ($signed(io_mulInput) * $signed(_14_25_inner_activation));
  assign _zz__zz__14_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_25_inner_macOut)) ? 16'h007f : _zz__14_25_inner_macOut_2);
  assign _zz__14_25_inner_macOut_2 = (($signed(_zz__14_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_25_inner_activation;
    end else begin
      io_macOut = _14_25_inner_macOut;
    end
  end

  assign _zz__14_25_inner_macOut = ($signed(_zz__zz__14_25_inner_macOut) + $signed(_zz__zz__14_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_25_inner_activation <= 8'h00;
      _14_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_25_inner_activation <= io_addInput;
      end else begin
        _14_25_inner_macOut <= _zz__14_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_472 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_24_inner_macOut;
  wire       [15:0]   _zz__zz__14_24_inner_macOut_1;
  wire       [15:0]   _zz__14_24_inner_macOut_1;
  wire       [15:0]   _zz__14_24_inner_macOut_2;
  reg        [7:0]    _14_24_inner_activation;
  reg        [7:0]    _14_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_24_inner_macOut;

  assign _zz__zz__14_24_inner_macOut = ($signed(io_mulInput) * $signed(_14_24_inner_activation));
  assign _zz__zz__14_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_24_inner_macOut)) ? 16'h007f : _zz__14_24_inner_macOut_2);
  assign _zz__14_24_inner_macOut_2 = (($signed(_zz__14_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_24_inner_activation;
    end else begin
      io_macOut = _14_24_inner_macOut;
    end
  end

  assign _zz__14_24_inner_macOut = ($signed(_zz__zz__14_24_inner_macOut) + $signed(_zz__zz__14_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_24_inner_activation <= 8'h00;
      _14_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_24_inner_activation <= io_addInput;
      end else begin
        _14_24_inner_macOut <= _zz__14_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_471 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_23_inner_macOut;
  wire       [15:0]   _zz__zz__14_23_inner_macOut_1;
  wire       [15:0]   _zz__14_23_inner_macOut_1;
  wire       [15:0]   _zz__14_23_inner_macOut_2;
  reg        [7:0]    _14_23_inner_activation;
  reg        [7:0]    _14_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_23_inner_macOut;

  assign _zz__zz__14_23_inner_macOut = ($signed(io_mulInput) * $signed(_14_23_inner_activation));
  assign _zz__zz__14_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_23_inner_macOut)) ? 16'h007f : _zz__14_23_inner_macOut_2);
  assign _zz__14_23_inner_macOut_2 = (($signed(_zz__14_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_23_inner_activation;
    end else begin
      io_macOut = _14_23_inner_macOut;
    end
  end

  assign _zz__14_23_inner_macOut = ($signed(_zz__zz__14_23_inner_macOut) + $signed(_zz__zz__14_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_23_inner_activation <= 8'h00;
      _14_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_23_inner_activation <= io_addInput;
      end else begin
        _14_23_inner_macOut <= _zz__14_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_470 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_22_inner_macOut;
  wire       [15:0]   _zz__zz__14_22_inner_macOut_1;
  wire       [15:0]   _zz__14_22_inner_macOut_1;
  wire       [15:0]   _zz__14_22_inner_macOut_2;
  reg        [7:0]    _14_22_inner_activation;
  reg        [7:0]    _14_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_22_inner_macOut;

  assign _zz__zz__14_22_inner_macOut = ($signed(io_mulInput) * $signed(_14_22_inner_activation));
  assign _zz__zz__14_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_22_inner_macOut)) ? 16'h007f : _zz__14_22_inner_macOut_2);
  assign _zz__14_22_inner_macOut_2 = (($signed(_zz__14_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_22_inner_activation;
    end else begin
      io_macOut = _14_22_inner_macOut;
    end
  end

  assign _zz__14_22_inner_macOut = ($signed(_zz__zz__14_22_inner_macOut) + $signed(_zz__zz__14_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_22_inner_activation <= 8'h00;
      _14_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_22_inner_activation <= io_addInput;
      end else begin
        _14_22_inner_macOut <= _zz__14_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_469 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_21_inner_macOut;
  wire       [15:0]   _zz__zz__14_21_inner_macOut_1;
  wire       [15:0]   _zz__14_21_inner_macOut_1;
  wire       [15:0]   _zz__14_21_inner_macOut_2;
  reg        [7:0]    _14_21_inner_activation;
  reg        [7:0]    _14_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_21_inner_macOut;

  assign _zz__zz__14_21_inner_macOut = ($signed(io_mulInput) * $signed(_14_21_inner_activation));
  assign _zz__zz__14_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_21_inner_macOut)) ? 16'h007f : _zz__14_21_inner_macOut_2);
  assign _zz__14_21_inner_macOut_2 = (($signed(_zz__14_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_21_inner_activation;
    end else begin
      io_macOut = _14_21_inner_macOut;
    end
  end

  assign _zz__14_21_inner_macOut = ($signed(_zz__zz__14_21_inner_macOut) + $signed(_zz__zz__14_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_21_inner_activation <= 8'h00;
      _14_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_21_inner_activation <= io_addInput;
      end else begin
        _14_21_inner_macOut <= _zz__14_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_468 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_20_inner_macOut;
  wire       [15:0]   _zz__zz__14_20_inner_macOut_1;
  wire       [15:0]   _zz__14_20_inner_macOut_1;
  wire       [15:0]   _zz__14_20_inner_macOut_2;
  reg        [7:0]    _14_20_inner_activation;
  reg        [7:0]    _14_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_20_inner_macOut;

  assign _zz__zz__14_20_inner_macOut = ($signed(io_mulInput) * $signed(_14_20_inner_activation));
  assign _zz__zz__14_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_20_inner_macOut)) ? 16'h007f : _zz__14_20_inner_macOut_2);
  assign _zz__14_20_inner_macOut_2 = (($signed(_zz__14_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_20_inner_activation;
    end else begin
      io_macOut = _14_20_inner_macOut;
    end
  end

  assign _zz__14_20_inner_macOut = ($signed(_zz__zz__14_20_inner_macOut) + $signed(_zz__zz__14_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_20_inner_activation <= 8'h00;
      _14_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_20_inner_activation <= io_addInput;
      end else begin
        _14_20_inner_macOut <= _zz__14_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_467 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_19_inner_macOut;
  wire       [15:0]   _zz__zz__14_19_inner_macOut_1;
  wire       [15:0]   _zz__14_19_inner_macOut_1;
  wire       [15:0]   _zz__14_19_inner_macOut_2;
  reg        [7:0]    _14_19_inner_activation;
  reg        [7:0]    _14_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_19_inner_macOut;

  assign _zz__zz__14_19_inner_macOut = ($signed(io_mulInput) * $signed(_14_19_inner_activation));
  assign _zz__zz__14_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_19_inner_macOut)) ? 16'h007f : _zz__14_19_inner_macOut_2);
  assign _zz__14_19_inner_macOut_2 = (($signed(_zz__14_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_19_inner_activation;
    end else begin
      io_macOut = _14_19_inner_macOut;
    end
  end

  assign _zz__14_19_inner_macOut = ($signed(_zz__zz__14_19_inner_macOut) + $signed(_zz__zz__14_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_19_inner_activation <= 8'h00;
      _14_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_19_inner_activation <= io_addInput;
      end else begin
        _14_19_inner_macOut <= _zz__14_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_466 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_18_inner_macOut;
  wire       [15:0]   _zz__zz__14_18_inner_macOut_1;
  wire       [15:0]   _zz__14_18_inner_macOut_1;
  wire       [15:0]   _zz__14_18_inner_macOut_2;
  reg        [7:0]    _14_18_inner_activation;
  reg        [7:0]    _14_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_18_inner_macOut;

  assign _zz__zz__14_18_inner_macOut = ($signed(io_mulInput) * $signed(_14_18_inner_activation));
  assign _zz__zz__14_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_18_inner_macOut)) ? 16'h007f : _zz__14_18_inner_macOut_2);
  assign _zz__14_18_inner_macOut_2 = (($signed(_zz__14_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_18_inner_activation;
    end else begin
      io_macOut = _14_18_inner_macOut;
    end
  end

  assign _zz__14_18_inner_macOut = ($signed(_zz__zz__14_18_inner_macOut) + $signed(_zz__zz__14_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_18_inner_activation <= 8'h00;
      _14_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_18_inner_activation <= io_addInput;
      end else begin
        _14_18_inner_macOut <= _zz__14_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_465 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_17_inner_macOut;
  wire       [15:0]   _zz__zz__14_17_inner_macOut_1;
  wire       [15:0]   _zz__14_17_inner_macOut_1;
  wire       [15:0]   _zz__14_17_inner_macOut_2;
  reg        [7:0]    _14_17_inner_activation;
  reg        [7:0]    _14_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_17_inner_macOut;

  assign _zz__zz__14_17_inner_macOut = ($signed(io_mulInput) * $signed(_14_17_inner_activation));
  assign _zz__zz__14_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_17_inner_macOut)) ? 16'h007f : _zz__14_17_inner_macOut_2);
  assign _zz__14_17_inner_macOut_2 = (($signed(_zz__14_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_17_inner_activation;
    end else begin
      io_macOut = _14_17_inner_macOut;
    end
  end

  assign _zz__14_17_inner_macOut = ($signed(_zz__zz__14_17_inner_macOut) + $signed(_zz__zz__14_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_17_inner_activation <= 8'h00;
      _14_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_17_inner_activation <= io_addInput;
      end else begin
        _14_17_inner_macOut <= _zz__14_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_464 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_16_inner_macOut;
  wire       [15:0]   _zz__zz__14_16_inner_macOut_1;
  wire       [15:0]   _zz__14_16_inner_macOut_1;
  wire       [15:0]   _zz__14_16_inner_macOut_2;
  reg        [7:0]    _14_16_inner_activation;
  reg        [7:0]    _14_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_16_inner_macOut;

  assign _zz__zz__14_16_inner_macOut = ($signed(io_mulInput) * $signed(_14_16_inner_activation));
  assign _zz__zz__14_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_16_inner_macOut)) ? 16'h007f : _zz__14_16_inner_macOut_2);
  assign _zz__14_16_inner_macOut_2 = (($signed(_zz__14_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_16_inner_activation;
    end else begin
      io_macOut = _14_16_inner_macOut;
    end
  end

  assign _zz__14_16_inner_macOut = ($signed(_zz__zz__14_16_inner_macOut) + $signed(_zz__zz__14_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_16_inner_activation <= 8'h00;
      _14_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_16_inner_activation <= io_addInput;
      end else begin
        _14_16_inner_macOut <= _zz__14_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_463 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_15_inner_macOut;
  wire       [15:0]   _zz__zz__14_15_inner_macOut_1;
  wire       [15:0]   _zz__14_15_inner_macOut_1;
  wire       [15:0]   _zz__14_15_inner_macOut_2;
  reg        [7:0]    _14_15_inner_activation;
  reg        [7:0]    _14_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_15_inner_macOut;

  assign _zz__zz__14_15_inner_macOut = ($signed(io_mulInput) * $signed(_14_15_inner_activation));
  assign _zz__zz__14_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_15_inner_macOut)) ? 16'h007f : _zz__14_15_inner_macOut_2);
  assign _zz__14_15_inner_macOut_2 = (($signed(_zz__14_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_15_inner_activation;
    end else begin
      io_macOut = _14_15_inner_macOut;
    end
  end

  assign _zz__14_15_inner_macOut = ($signed(_zz__zz__14_15_inner_macOut) + $signed(_zz__zz__14_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_15_inner_activation <= 8'h00;
      _14_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_15_inner_activation <= io_addInput;
      end else begin
        _14_15_inner_macOut <= _zz__14_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_462 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_14_inner_macOut;
  wire       [15:0]   _zz__zz__14_14_inner_macOut_1;
  wire       [15:0]   _zz__14_14_inner_macOut_1;
  wire       [15:0]   _zz__14_14_inner_macOut_2;
  reg        [7:0]    _14_14_inner_activation;
  reg        [7:0]    _14_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_14_inner_macOut;

  assign _zz__zz__14_14_inner_macOut = ($signed(io_mulInput) * $signed(_14_14_inner_activation));
  assign _zz__zz__14_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_14_inner_macOut)) ? 16'h007f : _zz__14_14_inner_macOut_2);
  assign _zz__14_14_inner_macOut_2 = (($signed(_zz__14_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_14_inner_activation;
    end else begin
      io_macOut = _14_14_inner_macOut;
    end
  end

  assign _zz__14_14_inner_macOut = ($signed(_zz__zz__14_14_inner_macOut) + $signed(_zz__zz__14_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_14_inner_activation <= 8'h00;
      _14_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_14_inner_activation <= io_addInput;
      end else begin
        _14_14_inner_macOut <= _zz__14_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_461 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_13_inner_macOut;
  wire       [15:0]   _zz__zz__14_13_inner_macOut_1;
  wire       [15:0]   _zz__14_13_inner_macOut_1;
  wire       [15:0]   _zz__14_13_inner_macOut_2;
  reg        [7:0]    _14_13_inner_activation;
  reg        [7:0]    _14_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_13_inner_macOut;

  assign _zz__zz__14_13_inner_macOut = ($signed(io_mulInput) * $signed(_14_13_inner_activation));
  assign _zz__zz__14_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_13_inner_macOut)) ? 16'h007f : _zz__14_13_inner_macOut_2);
  assign _zz__14_13_inner_macOut_2 = (($signed(_zz__14_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_13_inner_activation;
    end else begin
      io_macOut = _14_13_inner_macOut;
    end
  end

  assign _zz__14_13_inner_macOut = ($signed(_zz__zz__14_13_inner_macOut) + $signed(_zz__zz__14_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_13_inner_activation <= 8'h00;
      _14_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_13_inner_activation <= io_addInput;
      end else begin
        _14_13_inner_macOut <= _zz__14_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_460 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_12_inner_macOut;
  wire       [15:0]   _zz__zz__14_12_inner_macOut_1;
  wire       [15:0]   _zz__14_12_inner_macOut_1;
  wire       [15:0]   _zz__14_12_inner_macOut_2;
  reg        [7:0]    _14_12_inner_activation;
  reg        [7:0]    _14_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_12_inner_macOut;

  assign _zz__zz__14_12_inner_macOut = ($signed(io_mulInput) * $signed(_14_12_inner_activation));
  assign _zz__zz__14_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_12_inner_macOut)) ? 16'h007f : _zz__14_12_inner_macOut_2);
  assign _zz__14_12_inner_macOut_2 = (($signed(_zz__14_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_12_inner_activation;
    end else begin
      io_macOut = _14_12_inner_macOut;
    end
  end

  assign _zz__14_12_inner_macOut = ($signed(_zz__zz__14_12_inner_macOut) + $signed(_zz__zz__14_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_12_inner_activation <= 8'h00;
      _14_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_12_inner_activation <= io_addInput;
      end else begin
        _14_12_inner_macOut <= _zz__14_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_459 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_11_inner_macOut;
  wire       [15:0]   _zz__zz__14_11_inner_macOut_1;
  wire       [15:0]   _zz__14_11_inner_macOut_1;
  wire       [15:0]   _zz__14_11_inner_macOut_2;
  reg        [7:0]    _14_11_inner_activation;
  reg        [7:0]    _14_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_11_inner_macOut;

  assign _zz__zz__14_11_inner_macOut = ($signed(io_mulInput) * $signed(_14_11_inner_activation));
  assign _zz__zz__14_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_11_inner_macOut)) ? 16'h007f : _zz__14_11_inner_macOut_2);
  assign _zz__14_11_inner_macOut_2 = (($signed(_zz__14_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_11_inner_activation;
    end else begin
      io_macOut = _14_11_inner_macOut;
    end
  end

  assign _zz__14_11_inner_macOut = ($signed(_zz__zz__14_11_inner_macOut) + $signed(_zz__zz__14_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_11_inner_activation <= 8'h00;
      _14_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_11_inner_activation <= io_addInput;
      end else begin
        _14_11_inner_macOut <= _zz__14_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_458 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_10_inner_macOut;
  wire       [15:0]   _zz__zz__14_10_inner_macOut_1;
  wire       [15:0]   _zz__14_10_inner_macOut_1;
  wire       [15:0]   _zz__14_10_inner_macOut_2;
  reg        [7:0]    _14_10_inner_activation;
  reg        [7:0]    _14_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_10_inner_macOut;

  assign _zz__zz__14_10_inner_macOut = ($signed(io_mulInput) * $signed(_14_10_inner_activation));
  assign _zz__zz__14_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_10_inner_macOut)) ? 16'h007f : _zz__14_10_inner_macOut_2);
  assign _zz__14_10_inner_macOut_2 = (($signed(_zz__14_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_10_inner_activation;
    end else begin
      io_macOut = _14_10_inner_macOut;
    end
  end

  assign _zz__14_10_inner_macOut = ($signed(_zz__zz__14_10_inner_macOut) + $signed(_zz__zz__14_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_10_inner_activation <= 8'h00;
      _14_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_10_inner_activation <= io_addInput;
      end else begin
        _14_10_inner_macOut <= _zz__14_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_457 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_9_inner_macOut;
  wire       [15:0]   _zz__zz__14_9_inner_macOut_1;
  wire       [15:0]   _zz__14_9_inner_macOut_1;
  wire       [15:0]   _zz__14_9_inner_macOut_2;
  reg        [7:0]    _14_9_inner_activation;
  reg        [7:0]    _14_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_9_inner_macOut;

  assign _zz__zz__14_9_inner_macOut = ($signed(io_mulInput) * $signed(_14_9_inner_activation));
  assign _zz__zz__14_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_9_inner_macOut)) ? 16'h007f : _zz__14_9_inner_macOut_2);
  assign _zz__14_9_inner_macOut_2 = (($signed(_zz__14_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_9_inner_activation;
    end else begin
      io_macOut = _14_9_inner_macOut;
    end
  end

  assign _zz__14_9_inner_macOut = ($signed(_zz__zz__14_9_inner_macOut) + $signed(_zz__zz__14_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_9_inner_activation <= 8'h00;
      _14_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_9_inner_activation <= io_addInput;
      end else begin
        _14_9_inner_macOut <= _zz__14_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_456 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_8_inner_macOut;
  wire       [15:0]   _zz__zz__14_8_inner_macOut_1;
  wire       [15:0]   _zz__14_8_inner_macOut_1;
  wire       [15:0]   _zz__14_8_inner_macOut_2;
  reg        [7:0]    _14_8_inner_activation;
  reg        [7:0]    _14_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_8_inner_macOut;

  assign _zz__zz__14_8_inner_macOut = ($signed(io_mulInput) * $signed(_14_8_inner_activation));
  assign _zz__zz__14_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_8_inner_macOut)) ? 16'h007f : _zz__14_8_inner_macOut_2);
  assign _zz__14_8_inner_macOut_2 = (($signed(_zz__14_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_8_inner_activation;
    end else begin
      io_macOut = _14_8_inner_macOut;
    end
  end

  assign _zz__14_8_inner_macOut = ($signed(_zz__zz__14_8_inner_macOut) + $signed(_zz__zz__14_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_8_inner_activation <= 8'h00;
      _14_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_8_inner_activation <= io_addInput;
      end else begin
        _14_8_inner_macOut <= _zz__14_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_455 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_7_inner_macOut;
  wire       [15:0]   _zz__zz__14_7_inner_macOut_1;
  wire       [15:0]   _zz__14_7_inner_macOut_1;
  wire       [15:0]   _zz__14_7_inner_macOut_2;
  reg        [7:0]    _14_7_inner_activation;
  reg        [7:0]    _14_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_7_inner_macOut;

  assign _zz__zz__14_7_inner_macOut = ($signed(io_mulInput) * $signed(_14_7_inner_activation));
  assign _zz__zz__14_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_7_inner_macOut)) ? 16'h007f : _zz__14_7_inner_macOut_2);
  assign _zz__14_7_inner_macOut_2 = (($signed(_zz__14_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_7_inner_activation;
    end else begin
      io_macOut = _14_7_inner_macOut;
    end
  end

  assign _zz__14_7_inner_macOut = ($signed(_zz__zz__14_7_inner_macOut) + $signed(_zz__zz__14_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_7_inner_activation <= 8'h00;
      _14_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_7_inner_activation <= io_addInput;
      end else begin
        _14_7_inner_macOut <= _zz__14_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_454 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_6_inner_macOut;
  wire       [15:0]   _zz__zz__14_6_inner_macOut_1;
  wire       [15:0]   _zz__14_6_inner_macOut_1;
  wire       [15:0]   _zz__14_6_inner_macOut_2;
  reg        [7:0]    _14_6_inner_activation;
  reg        [7:0]    _14_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_6_inner_macOut;

  assign _zz__zz__14_6_inner_macOut = ($signed(io_mulInput) * $signed(_14_6_inner_activation));
  assign _zz__zz__14_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_6_inner_macOut)) ? 16'h007f : _zz__14_6_inner_macOut_2);
  assign _zz__14_6_inner_macOut_2 = (($signed(_zz__14_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_6_inner_activation;
    end else begin
      io_macOut = _14_6_inner_macOut;
    end
  end

  assign _zz__14_6_inner_macOut = ($signed(_zz__zz__14_6_inner_macOut) + $signed(_zz__zz__14_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_6_inner_activation <= 8'h00;
      _14_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_6_inner_activation <= io_addInput;
      end else begin
        _14_6_inner_macOut <= _zz__14_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_453 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_5_inner_macOut;
  wire       [15:0]   _zz__zz__14_5_inner_macOut_1;
  wire       [15:0]   _zz__14_5_inner_macOut_1;
  wire       [15:0]   _zz__14_5_inner_macOut_2;
  reg        [7:0]    _14_5_inner_activation;
  reg        [7:0]    _14_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_5_inner_macOut;

  assign _zz__zz__14_5_inner_macOut = ($signed(io_mulInput) * $signed(_14_5_inner_activation));
  assign _zz__zz__14_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_5_inner_macOut)) ? 16'h007f : _zz__14_5_inner_macOut_2);
  assign _zz__14_5_inner_macOut_2 = (($signed(_zz__14_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_5_inner_activation;
    end else begin
      io_macOut = _14_5_inner_macOut;
    end
  end

  assign _zz__14_5_inner_macOut = ($signed(_zz__zz__14_5_inner_macOut) + $signed(_zz__zz__14_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_5_inner_activation <= 8'h00;
      _14_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_5_inner_activation <= io_addInput;
      end else begin
        _14_5_inner_macOut <= _zz__14_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_452 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_4_inner_macOut;
  wire       [15:0]   _zz__zz__14_4_inner_macOut_1;
  wire       [15:0]   _zz__14_4_inner_macOut_1;
  wire       [15:0]   _zz__14_4_inner_macOut_2;
  reg        [7:0]    _14_4_inner_activation;
  reg        [7:0]    _14_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_4_inner_macOut;

  assign _zz__zz__14_4_inner_macOut = ($signed(io_mulInput) * $signed(_14_4_inner_activation));
  assign _zz__zz__14_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_4_inner_macOut)) ? 16'h007f : _zz__14_4_inner_macOut_2);
  assign _zz__14_4_inner_macOut_2 = (($signed(_zz__14_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_4_inner_activation;
    end else begin
      io_macOut = _14_4_inner_macOut;
    end
  end

  assign _zz__14_4_inner_macOut = ($signed(_zz__zz__14_4_inner_macOut) + $signed(_zz__zz__14_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_4_inner_activation <= 8'h00;
      _14_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_4_inner_activation <= io_addInput;
      end else begin
        _14_4_inner_macOut <= _zz__14_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_451 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_3_inner_macOut;
  wire       [15:0]   _zz__zz__14_3_inner_macOut_1;
  wire       [15:0]   _zz__14_3_inner_macOut_1;
  wire       [15:0]   _zz__14_3_inner_macOut_2;
  reg        [7:0]    _14_3_inner_activation;
  reg        [7:0]    _14_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_3_inner_macOut;

  assign _zz__zz__14_3_inner_macOut = ($signed(io_mulInput) * $signed(_14_3_inner_activation));
  assign _zz__zz__14_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_3_inner_macOut)) ? 16'h007f : _zz__14_3_inner_macOut_2);
  assign _zz__14_3_inner_macOut_2 = (($signed(_zz__14_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_3_inner_activation;
    end else begin
      io_macOut = _14_3_inner_macOut;
    end
  end

  assign _zz__14_3_inner_macOut = ($signed(_zz__zz__14_3_inner_macOut) + $signed(_zz__zz__14_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_3_inner_activation <= 8'h00;
      _14_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_3_inner_activation <= io_addInput;
      end else begin
        _14_3_inner_macOut <= _zz__14_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_450 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_2_inner_macOut;
  wire       [15:0]   _zz__zz__14_2_inner_macOut_1;
  wire       [15:0]   _zz__14_2_inner_macOut_1;
  wire       [15:0]   _zz__14_2_inner_macOut_2;
  reg        [7:0]    _14_2_inner_activation;
  reg        [7:0]    _14_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_2_inner_macOut;

  assign _zz__zz__14_2_inner_macOut = ($signed(io_mulInput) * $signed(_14_2_inner_activation));
  assign _zz__zz__14_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_2_inner_macOut)) ? 16'h007f : _zz__14_2_inner_macOut_2);
  assign _zz__14_2_inner_macOut_2 = (($signed(_zz__14_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_2_inner_activation;
    end else begin
      io_macOut = _14_2_inner_macOut;
    end
  end

  assign _zz__14_2_inner_macOut = ($signed(_zz__zz__14_2_inner_macOut) + $signed(_zz__zz__14_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_2_inner_activation <= 8'h00;
      _14_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_2_inner_activation <= io_addInput;
      end else begin
        _14_2_inner_macOut <= _zz__14_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_449 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_1_inner_macOut;
  wire       [15:0]   _zz__zz__14_1_inner_macOut_1;
  wire       [15:0]   _zz__14_1_inner_macOut_1;
  wire       [15:0]   _zz__14_1_inner_macOut_2;
  reg        [7:0]    _14_1_inner_activation;
  reg        [7:0]    _14_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_1_inner_macOut;

  assign _zz__zz__14_1_inner_macOut = ($signed(io_mulInput) * $signed(_14_1_inner_activation));
  assign _zz__zz__14_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_1_inner_macOut)) ? 16'h007f : _zz__14_1_inner_macOut_2);
  assign _zz__14_1_inner_macOut_2 = (($signed(_zz__14_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_1_inner_activation;
    end else begin
      io_macOut = _14_1_inner_macOut;
    end
  end

  assign _zz__14_1_inner_macOut = ($signed(_zz__zz__14_1_inner_macOut) + $signed(_zz__zz__14_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_1_inner_activation <= 8'h00;
      _14_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_1_inner_activation <= io_addInput;
      end else begin
        _14_1_inner_macOut <= _zz__14_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_448 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__14_0_inner_macOut;
  wire       [15:0]   _zz__zz__14_0_inner_macOut_1;
  wire       [15:0]   _zz__14_0_inner_macOut_1;
  wire       [15:0]   _zz__14_0_inner_macOut_2;
  reg        [7:0]    _14_0_inner_activation;
  reg        [7:0]    _14_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__14_0_inner_macOut;

  assign _zz__zz__14_0_inner_macOut = ($signed(io_mulInput) * $signed(_14_0_inner_activation));
  assign _zz__zz__14_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__14_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__14_0_inner_macOut)) ? 16'h007f : _zz__14_0_inner_macOut_2);
  assign _zz__14_0_inner_macOut_2 = (($signed(_zz__14_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__14_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _14_0_inner_activation;
    end else begin
      io_macOut = _14_0_inner_macOut;
    end
  end

  assign _zz__14_0_inner_macOut = ($signed(_zz__zz__14_0_inner_macOut) + $signed(_zz__zz__14_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _14_0_inner_activation <= 8'h00;
      _14_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _14_0_inner_activation <= io_addInput;
      end else begin
        _14_0_inner_macOut <= _zz__14_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_447 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_31_inner_macOut;
  wire       [15:0]   _zz__zz__13_31_inner_macOut_1;
  wire       [15:0]   _zz__13_31_inner_macOut_1;
  wire       [15:0]   _zz__13_31_inner_macOut_2;
  reg        [7:0]    _13_31_inner_activation;
  reg        [7:0]    _13_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_31_inner_macOut;

  assign _zz__zz__13_31_inner_macOut = ($signed(io_mulInput) * $signed(_13_31_inner_activation));
  assign _zz__zz__13_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_31_inner_macOut)) ? 16'h007f : _zz__13_31_inner_macOut_2);
  assign _zz__13_31_inner_macOut_2 = (($signed(_zz__13_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_31_inner_activation;
    end else begin
      io_macOut = _13_31_inner_macOut;
    end
  end

  assign _zz__13_31_inner_macOut = ($signed(_zz__zz__13_31_inner_macOut) + $signed(_zz__zz__13_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_31_inner_activation <= 8'h00;
      _13_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_31_inner_activation <= io_addInput;
      end else begin
        _13_31_inner_macOut <= _zz__13_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_446 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_30_inner_macOut;
  wire       [15:0]   _zz__zz__13_30_inner_macOut_1;
  wire       [15:0]   _zz__13_30_inner_macOut_1;
  wire       [15:0]   _zz__13_30_inner_macOut_2;
  reg        [7:0]    _13_30_inner_activation;
  reg        [7:0]    _13_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_30_inner_macOut;

  assign _zz__zz__13_30_inner_macOut = ($signed(io_mulInput) * $signed(_13_30_inner_activation));
  assign _zz__zz__13_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_30_inner_macOut)) ? 16'h007f : _zz__13_30_inner_macOut_2);
  assign _zz__13_30_inner_macOut_2 = (($signed(_zz__13_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_30_inner_activation;
    end else begin
      io_macOut = _13_30_inner_macOut;
    end
  end

  assign _zz__13_30_inner_macOut = ($signed(_zz__zz__13_30_inner_macOut) + $signed(_zz__zz__13_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_30_inner_activation <= 8'h00;
      _13_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_30_inner_activation <= io_addInput;
      end else begin
        _13_30_inner_macOut <= _zz__13_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_445 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_29_inner_macOut;
  wire       [15:0]   _zz__zz__13_29_inner_macOut_1;
  wire       [15:0]   _zz__13_29_inner_macOut_1;
  wire       [15:0]   _zz__13_29_inner_macOut_2;
  reg        [7:0]    _13_29_inner_activation;
  reg        [7:0]    _13_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_29_inner_macOut;

  assign _zz__zz__13_29_inner_macOut = ($signed(io_mulInput) * $signed(_13_29_inner_activation));
  assign _zz__zz__13_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_29_inner_macOut)) ? 16'h007f : _zz__13_29_inner_macOut_2);
  assign _zz__13_29_inner_macOut_2 = (($signed(_zz__13_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_29_inner_activation;
    end else begin
      io_macOut = _13_29_inner_macOut;
    end
  end

  assign _zz__13_29_inner_macOut = ($signed(_zz__zz__13_29_inner_macOut) + $signed(_zz__zz__13_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_29_inner_activation <= 8'h00;
      _13_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_29_inner_activation <= io_addInput;
      end else begin
        _13_29_inner_macOut <= _zz__13_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_444 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_28_inner_macOut;
  wire       [15:0]   _zz__zz__13_28_inner_macOut_1;
  wire       [15:0]   _zz__13_28_inner_macOut_1;
  wire       [15:0]   _zz__13_28_inner_macOut_2;
  reg        [7:0]    _13_28_inner_activation;
  reg        [7:0]    _13_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_28_inner_macOut;

  assign _zz__zz__13_28_inner_macOut = ($signed(io_mulInput) * $signed(_13_28_inner_activation));
  assign _zz__zz__13_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_28_inner_macOut)) ? 16'h007f : _zz__13_28_inner_macOut_2);
  assign _zz__13_28_inner_macOut_2 = (($signed(_zz__13_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_28_inner_activation;
    end else begin
      io_macOut = _13_28_inner_macOut;
    end
  end

  assign _zz__13_28_inner_macOut = ($signed(_zz__zz__13_28_inner_macOut) + $signed(_zz__zz__13_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_28_inner_activation <= 8'h00;
      _13_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_28_inner_activation <= io_addInput;
      end else begin
        _13_28_inner_macOut <= _zz__13_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_443 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_27_inner_macOut;
  wire       [15:0]   _zz__zz__13_27_inner_macOut_1;
  wire       [15:0]   _zz__13_27_inner_macOut_1;
  wire       [15:0]   _zz__13_27_inner_macOut_2;
  reg        [7:0]    _13_27_inner_activation;
  reg        [7:0]    _13_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_27_inner_macOut;

  assign _zz__zz__13_27_inner_macOut = ($signed(io_mulInput) * $signed(_13_27_inner_activation));
  assign _zz__zz__13_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_27_inner_macOut)) ? 16'h007f : _zz__13_27_inner_macOut_2);
  assign _zz__13_27_inner_macOut_2 = (($signed(_zz__13_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_27_inner_activation;
    end else begin
      io_macOut = _13_27_inner_macOut;
    end
  end

  assign _zz__13_27_inner_macOut = ($signed(_zz__zz__13_27_inner_macOut) + $signed(_zz__zz__13_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_27_inner_activation <= 8'h00;
      _13_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_27_inner_activation <= io_addInput;
      end else begin
        _13_27_inner_macOut <= _zz__13_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_442 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_26_inner_macOut;
  wire       [15:0]   _zz__zz__13_26_inner_macOut_1;
  wire       [15:0]   _zz__13_26_inner_macOut_1;
  wire       [15:0]   _zz__13_26_inner_macOut_2;
  reg        [7:0]    _13_26_inner_activation;
  reg        [7:0]    _13_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_26_inner_macOut;

  assign _zz__zz__13_26_inner_macOut = ($signed(io_mulInput) * $signed(_13_26_inner_activation));
  assign _zz__zz__13_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_26_inner_macOut)) ? 16'h007f : _zz__13_26_inner_macOut_2);
  assign _zz__13_26_inner_macOut_2 = (($signed(_zz__13_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_26_inner_activation;
    end else begin
      io_macOut = _13_26_inner_macOut;
    end
  end

  assign _zz__13_26_inner_macOut = ($signed(_zz__zz__13_26_inner_macOut) + $signed(_zz__zz__13_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_26_inner_activation <= 8'h00;
      _13_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_26_inner_activation <= io_addInput;
      end else begin
        _13_26_inner_macOut <= _zz__13_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_441 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_25_inner_macOut;
  wire       [15:0]   _zz__zz__13_25_inner_macOut_1;
  wire       [15:0]   _zz__13_25_inner_macOut_1;
  wire       [15:0]   _zz__13_25_inner_macOut_2;
  reg        [7:0]    _13_25_inner_activation;
  reg        [7:0]    _13_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_25_inner_macOut;

  assign _zz__zz__13_25_inner_macOut = ($signed(io_mulInput) * $signed(_13_25_inner_activation));
  assign _zz__zz__13_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_25_inner_macOut)) ? 16'h007f : _zz__13_25_inner_macOut_2);
  assign _zz__13_25_inner_macOut_2 = (($signed(_zz__13_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_25_inner_activation;
    end else begin
      io_macOut = _13_25_inner_macOut;
    end
  end

  assign _zz__13_25_inner_macOut = ($signed(_zz__zz__13_25_inner_macOut) + $signed(_zz__zz__13_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_25_inner_activation <= 8'h00;
      _13_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_25_inner_activation <= io_addInput;
      end else begin
        _13_25_inner_macOut <= _zz__13_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_440 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_24_inner_macOut;
  wire       [15:0]   _zz__zz__13_24_inner_macOut_1;
  wire       [15:0]   _zz__13_24_inner_macOut_1;
  wire       [15:0]   _zz__13_24_inner_macOut_2;
  reg        [7:0]    _13_24_inner_activation;
  reg        [7:0]    _13_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_24_inner_macOut;

  assign _zz__zz__13_24_inner_macOut = ($signed(io_mulInput) * $signed(_13_24_inner_activation));
  assign _zz__zz__13_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_24_inner_macOut)) ? 16'h007f : _zz__13_24_inner_macOut_2);
  assign _zz__13_24_inner_macOut_2 = (($signed(_zz__13_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_24_inner_activation;
    end else begin
      io_macOut = _13_24_inner_macOut;
    end
  end

  assign _zz__13_24_inner_macOut = ($signed(_zz__zz__13_24_inner_macOut) + $signed(_zz__zz__13_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_24_inner_activation <= 8'h00;
      _13_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_24_inner_activation <= io_addInput;
      end else begin
        _13_24_inner_macOut <= _zz__13_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_439 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_23_inner_macOut;
  wire       [15:0]   _zz__zz__13_23_inner_macOut_1;
  wire       [15:0]   _zz__13_23_inner_macOut_1;
  wire       [15:0]   _zz__13_23_inner_macOut_2;
  reg        [7:0]    _13_23_inner_activation;
  reg        [7:0]    _13_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_23_inner_macOut;

  assign _zz__zz__13_23_inner_macOut = ($signed(io_mulInput) * $signed(_13_23_inner_activation));
  assign _zz__zz__13_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_23_inner_macOut)) ? 16'h007f : _zz__13_23_inner_macOut_2);
  assign _zz__13_23_inner_macOut_2 = (($signed(_zz__13_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_23_inner_activation;
    end else begin
      io_macOut = _13_23_inner_macOut;
    end
  end

  assign _zz__13_23_inner_macOut = ($signed(_zz__zz__13_23_inner_macOut) + $signed(_zz__zz__13_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_23_inner_activation <= 8'h00;
      _13_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_23_inner_activation <= io_addInput;
      end else begin
        _13_23_inner_macOut <= _zz__13_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_438 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_22_inner_macOut;
  wire       [15:0]   _zz__zz__13_22_inner_macOut_1;
  wire       [15:0]   _zz__13_22_inner_macOut_1;
  wire       [15:0]   _zz__13_22_inner_macOut_2;
  reg        [7:0]    _13_22_inner_activation;
  reg        [7:0]    _13_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_22_inner_macOut;

  assign _zz__zz__13_22_inner_macOut = ($signed(io_mulInput) * $signed(_13_22_inner_activation));
  assign _zz__zz__13_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_22_inner_macOut)) ? 16'h007f : _zz__13_22_inner_macOut_2);
  assign _zz__13_22_inner_macOut_2 = (($signed(_zz__13_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_22_inner_activation;
    end else begin
      io_macOut = _13_22_inner_macOut;
    end
  end

  assign _zz__13_22_inner_macOut = ($signed(_zz__zz__13_22_inner_macOut) + $signed(_zz__zz__13_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_22_inner_activation <= 8'h00;
      _13_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_22_inner_activation <= io_addInput;
      end else begin
        _13_22_inner_macOut <= _zz__13_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_437 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_21_inner_macOut;
  wire       [15:0]   _zz__zz__13_21_inner_macOut_1;
  wire       [15:0]   _zz__13_21_inner_macOut_1;
  wire       [15:0]   _zz__13_21_inner_macOut_2;
  reg        [7:0]    _13_21_inner_activation;
  reg        [7:0]    _13_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_21_inner_macOut;

  assign _zz__zz__13_21_inner_macOut = ($signed(io_mulInput) * $signed(_13_21_inner_activation));
  assign _zz__zz__13_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_21_inner_macOut)) ? 16'h007f : _zz__13_21_inner_macOut_2);
  assign _zz__13_21_inner_macOut_2 = (($signed(_zz__13_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_21_inner_activation;
    end else begin
      io_macOut = _13_21_inner_macOut;
    end
  end

  assign _zz__13_21_inner_macOut = ($signed(_zz__zz__13_21_inner_macOut) + $signed(_zz__zz__13_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_21_inner_activation <= 8'h00;
      _13_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_21_inner_activation <= io_addInput;
      end else begin
        _13_21_inner_macOut <= _zz__13_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_436 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_20_inner_macOut;
  wire       [15:0]   _zz__zz__13_20_inner_macOut_1;
  wire       [15:0]   _zz__13_20_inner_macOut_1;
  wire       [15:0]   _zz__13_20_inner_macOut_2;
  reg        [7:0]    _13_20_inner_activation;
  reg        [7:0]    _13_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_20_inner_macOut;

  assign _zz__zz__13_20_inner_macOut = ($signed(io_mulInput) * $signed(_13_20_inner_activation));
  assign _zz__zz__13_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_20_inner_macOut)) ? 16'h007f : _zz__13_20_inner_macOut_2);
  assign _zz__13_20_inner_macOut_2 = (($signed(_zz__13_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_20_inner_activation;
    end else begin
      io_macOut = _13_20_inner_macOut;
    end
  end

  assign _zz__13_20_inner_macOut = ($signed(_zz__zz__13_20_inner_macOut) + $signed(_zz__zz__13_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_20_inner_activation <= 8'h00;
      _13_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_20_inner_activation <= io_addInput;
      end else begin
        _13_20_inner_macOut <= _zz__13_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_435 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_19_inner_macOut;
  wire       [15:0]   _zz__zz__13_19_inner_macOut_1;
  wire       [15:0]   _zz__13_19_inner_macOut_1;
  wire       [15:0]   _zz__13_19_inner_macOut_2;
  reg        [7:0]    _13_19_inner_activation;
  reg        [7:0]    _13_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_19_inner_macOut;

  assign _zz__zz__13_19_inner_macOut = ($signed(io_mulInput) * $signed(_13_19_inner_activation));
  assign _zz__zz__13_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_19_inner_macOut)) ? 16'h007f : _zz__13_19_inner_macOut_2);
  assign _zz__13_19_inner_macOut_2 = (($signed(_zz__13_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_19_inner_activation;
    end else begin
      io_macOut = _13_19_inner_macOut;
    end
  end

  assign _zz__13_19_inner_macOut = ($signed(_zz__zz__13_19_inner_macOut) + $signed(_zz__zz__13_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_19_inner_activation <= 8'h00;
      _13_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_19_inner_activation <= io_addInput;
      end else begin
        _13_19_inner_macOut <= _zz__13_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_434 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_18_inner_macOut;
  wire       [15:0]   _zz__zz__13_18_inner_macOut_1;
  wire       [15:0]   _zz__13_18_inner_macOut_1;
  wire       [15:0]   _zz__13_18_inner_macOut_2;
  reg        [7:0]    _13_18_inner_activation;
  reg        [7:0]    _13_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_18_inner_macOut;

  assign _zz__zz__13_18_inner_macOut = ($signed(io_mulInput) * $signed(_13_18_inner_activation));
  assign _zz__zz__13_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_18_inner_macOut)) ? 16'h007f : _zz__13_18_inner_macOut_2);
  assign _zz__13_18_inner_macOut_2 = (($signed(_zz__13_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_18_inner_activation;
    end else begin
      io_macOut = _13_18_inner_macOut;
    end
  end

  assign _zz__13_18_inner_macOut = ($signed(_zz__zz__13_18_inner_macOut) + $signed(_zz__zz__13_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_18_inner_activation <= 8'h00;
      _13_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_18_inner_activation <= io_addInput;
      end else begin
        _13_18_inner_macOut <= _zz__13_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_433 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_17_inner_macOut;
  wire       [15:0]   _zz__zz__13_17_inner_macOut_1;
  wire       [15:0]   _zz__13_17_inner_macOut_1;
  wire       [15:0]   _zz__13_17_inner_macOut_2;
  reg        [7:0]    _13_17_inner_activation;
  reg        [7:0]    _13_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_17_inner_macOut;

  assign _zz__zz__13_17_inner_macOut = ($signed(io_mulInput) * $signed(_13_17_inner_activation));
  assign _zz__zz__13_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_17_inner_macOut)) ? 16'h007f : _zz__13_17_inner_macOut_2);
  assign _zz__13_17_inner_macOut_2 = (($signed(_zz__13_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_17_inner_activation;
    end else begin
      io_macOut = _13_17_inner_macOut;
    end
  end

  assign _zz__13_17_inner_macOut = ($signed(_zz__zz__13_17_inner_macOut) + $signed(_zz__zz__13_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_17_inner_activation <= 8'h00;
      _13_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_17_inner_activation <= io_addInput;
      end else begin
        _13_17_inner_macOut <= _zz__13_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_432 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_16_inner_macOut;
  wire       [15:0]   _zz__zz__13_16_inner_macOut_1;
  wire       [15:0]   _zz__13_16_inner_macOut_1;
  wire       [15:0]   _zz__13_16_inner_macOut_2;
  reg        [7:0]    _13_16_inner_activation;
  reg        [7:0]    _13_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_16_inner_macOut;

  assign _zz__zz__13_16_inner_macOut = ($signed(io_mulInput) * $signed(_13_16_inner_activation));
  assign _zz__zz__13_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_16_inner_macOut)) ? 16'h007f : _zz__13_16_inner_macOut_2);
  assign _zz__13_16_inner_macOut_2 = (($signed(_zz__13_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_16_inner_activation;
    end else begin
      io_macOut = _13_16_inner_macOut;
    end
  end

  assign _zz__13_16_inner_macOut = ($signed(_zz__zz__13_16_inner_macOut) + $signed(_zz__zz__13_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_16_inner_activation <= 8'h00;
      _13_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_16_inner_activation <= io_addInput;
      end else begin
        _13_16_inner_macOut <= _zz__13_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_431 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_15_inner_macOut;
  wire       [15:0]   _zz__zz__13_15_inner_macOut_1;
  wire       [15:0]   _zz__13_15_inner_macOut_1;
  wire       [15:0]   _zz__13_15_inner_macOut_2;
  reg        [7:0]    _13_15_inner_activation;
  reg        [7:0]    _13_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_15_inner_macOut;

  assign _zz__zz__13_15_inner_macOut = ($signed(io_mulInput) * $signed(_13_15_inner_activation));
  assign _zz__zz__13_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_15_inner_macOut)) ? 16'h007f : _zz__13_15_inner_macOut_2);
  assign _zz__13_15_inner_macOut_2 = (($signed(_zz__13_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_15_inner_activation;
    end else begin
      io_macOut = _13_15_inner_macOut;
    end
  end

  assign _zz__13_15_inner_macOut = ($signed(_zz__zz__13_15_inner_macOut) + $signed(_zz__zz__13_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_15_inner_activation <= 8'h00;
      _13_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_15_inner_activation <= io_addInput;
      end else begin
        _13_15_inner_macOut <= _zz__13_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_430 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_14_inner_macOut;
  wire       [15:0]   _zz__zz__13_14_inner_macOut_1;
  wire       [15:0]   _zz__13_14_inner_macOut_1;
  wire       [15:0]   _zz__13_14_inner_macOut_2;
  reg        [7:0]    _13_14_inner_activation;
  reg        [7:0]    _13_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_14_inner_macOut;

  assign _zz__zz__13_14_inner_macOut = ($signed(io_mulInput) * $signed(_13_14_inner_activation));
  assign _zz__zz__13_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_14_inner_macOut)) ? 16'h007f : _zz__13_14_inner_macOut_2);
  assign _zz__13_14_inner_macOut_2 = (($signed(_zz__13_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_14_inner_activation;
    end else begin
      io_macOut = _13_14_inner_macOut;
    end
  end

  assign _zz__13_14_inner_macOut = ($signed(_zz__zz__13_14_inner_macOut) + $signed(_zz__zz__13_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_14_inner_activation <= 8'h00;
      _13_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_14_inner_activation <= io_addInput;
      end else begin
        _13_14_inner_macOut <= _zz__13_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_429 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_13_inner_macOut;
  wire       [15:0]   _zz__zz__13_13_inner_macOut_1;
  wire       [15:0]   _zz__13_13_inner_macOut_1;
  wire       [15:0]   _zz__13_13_inner_macOut_2;
  reg        [7:0]    _13_13_inner_activation;
  reg        [7:0]    _13_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_13_inner_macOut;

  assign _zz__zz__13_13_inner_macOut = ($signed(io_mulInput) * $signed(_13_13_inner_activation));
  assign _zz__zz__13_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_13_inner_macOut)) ? 16'h007f : _zz__13_13_inner_macOut_2);
  assign _zz__13_13_inner_macOut_2 = (($signed(_zz__13_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_13_inner_activation;
    end else begin
      io_macOut = _13_13_inner_macOut;
    end
  end

  assign _zz__13_13_inner_macOut = ($signed(_zz__zz__13_13_inner_macOut) + $signed(_zz__zz__13_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_13_inner_activation <= 8'h00;
      _13_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_13_inner_activation <= io_addInput;
      end else begin
        _13_13_inner_macOut <= _zz__13_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_428 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_12_inner_macOut;
  wire       [15:0]   _zz__zz__13_12_inner_macOut_1;
  wire       [15:0]   _zz__13_12_inner_macOut_1;
  wire       [15:0]   _zz__13_12_inner_macOut_2;
  reg        [7:0]    _13_12_inner_activation;
  reg        [7:0]    _13_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_12_inner_macOut;

  assign _zz__zz__13_12_inner_macOut = ($signed(io_mulInput) * $signed(_13_12_inner_activation));
  assign _zz__zz__13_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_12_inner_macOut)) ? 16'h007f : _zz__13_12_inner_macOut_2);
  assign _zz__13_12_inner_macOut_2 = (($signed(_zz__13_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_12_inner_activation;
    end else begin
      io_macOut = _13_12_inner_macOut;
    end
  end

  assign _zz__13_12_inner_macOut = ($signed(_zz__zz__13_12_inner_macOut) + $signed(_zz__zz__13_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_12_inner_activation <= 8'h00;
      _13_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_12_inner_activation <= io_addInput;
      end else begin
        _13_12_inner_macOut <= _zz__13_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_427 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_11_inner_macOut;
  wire       [15:0]   _zz__zz__13_11_inner_macOut_1;
  wire       [15:0]   _zz__13_11_inner_macOut_1;
  wire       [15:0]   _zz__13_11_inner_macOut_2;
  reg        [7:0]    _13_11_inner_activation;
  reg        [7:0]    _13_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_11_inner_macOut;

  assign _zz__zz__13_11_inner_macOut = ($signed(io_mulInput) * $signed(_13_11_inner_activation));
  assign _zz__zz__13_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_11_inner_macOut)) ? 16'h007f : _zz__13_11_inner_macOut_2);
  assign _zz__13_11_inner_macOut_2 = (($signed(_zz__13_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_11_inner_activation;
    end else begin
      io_macOut = _13_11_inner_macOut;
    end
  end

  assign _zz__13_11_inner_macOut = ($signed(_zz__zz__13_11_inner_macOut) + $signed(_zz__zz__13_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_11_inner_activation <= 8'h00;
      _13_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_11_inner_activation <= io_addInput;
      end else begin
        _13_11_inner_macOut <= _zz__13_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_426 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_10_inner_macOut;
  wire       [15:0]   _zz__zz__13_10_inner_macOut_1;
  wire       [15:0]   _zz__13_10_inner_macOut_1;
  wire       [15:0]   _zz__13_10_inner_macOut_2;
  reg        [7:0]    _13_10_inner_activation;
  reg        [7:0]    _13_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_10_inner_macOut;

  assign _zz__zz__13_10_inner_macOut = ($signed(io_mulInput) * $signed(_13_10_inner_activation));
  assign _zz__zz__13_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_10_inner_macOut)) ? 16'h007f : _zz__13_10_inner_macOut_2);
  assign _zz__13_10_inner_macOut_2 = (($signed(_zz__13_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_10_inner_activation;
    end else begin
      io_macOut = _13_10_inner_macOut;
    end
  end

  assign _zz__13_10_inner_macOut = ($signed(_zz__zz__13_10_inner_macOut) + $signed(_zz__zz__13_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_10_inner_activation <= 8'h00;
      _13_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_10_inner_activation <= io_addInput;
      end else begin
        _13_10_inner_macOut <= _zz__13_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_425 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_9_inner_macOut;
  wire       [15:0]   _zz__zz__13_9_inner_macOut_1;
  wire       [15:0]   _zz__13_9_inner_macOut_1;
  wire       [15:0]   _zz__13_9_inner_macOut_2;
  reg        [7:0]    _13_9_inner_activation;
  reg        [7:0]    _13_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_9_inner_macOut;

  assign _zz__zz__13_9_inner_macOut = ($signed(io_mulInput) * $signed(_13_9_inner_activation));
  assign _zz__zz__13_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_9_inner_macOut)) ? 16'h007f : _zz__13_9_inner_macOut_2);
  assign _zz__13_9_inner_macOut_2 = (($signed(_zz__13_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_9_inner_activation;
    end else begin
      io_macOut = _13_9_inner_macOut;
    end
  end

  assign _zz__13_9_inner_macOut = ($signed(_zz__zz__13_9_inner_macOut) + $signed(_zz__zz__13_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_9_inner_activation <= 8'h00;
      _13_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_9_inner_activation <= io_addInput;
      end else begin
        _13_9_inner_macOut <= _zz__13_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_424 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_8_inner_macOut;
  wire       [15:0]   _zz__zz__13_8_inner_macOut_1;
  wire       [15:0]   _zz__13_8_inner_macOut_1;
  wire       [15:0]   _zz__13_8_inner_macOut_2;
  reg        [7:0]    _13_8_inner_activation;
  reg        [7:0]    _13_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_8_inner_macOut;

  assign _zz__zz__13_8_inner_macOut = ($signed(io_mulInput) * $signed(_13_8_inner_activation));
  assign _zz__zz__13_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_8_inner_macOut)) ? 16'h007f : _zz__13_8_inner_macOut_2);
  assign _zz__13_8_inner_macOut_2 = (($signed(_zz__13_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_8_inner_activation;
    end else begin
      io_macOut = _13_8_inner_macOut;
    end
  end

  assign _zz__13_8_inner_macOut = ($signed(_zz__zz__13_8_inner_macOut) + $signed(_zz__zz__13_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_8_inner_activation <= 8'h00;
      _13_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_8_inner_activation <= io_addInput;
      end else begin
        _13_8_inner_macOut <= _zz__13_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_423 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_7_inner_macOut;
  wire       [15:0]   _zz__zz__13_7_inner_macOut_1;
  wire       [15:0]   _zz__13_7_inner_macOut_1;
  wire       [15:0]   _zz__13_7_inner_macOut_2;
  reg        [7:0]    _13_7_inner_activation;
  reg        [7:0]    _13_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_7_inner_macOut;

  assign _zz__zz__13_7_inner_macOut = ($signed(io_mulInput) * $signed(_13_7_inner_activation));
  assign _zz__zz__13_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_7_inner_macOut)) ? 16'h007f : _zz__13_7_inner_macOut_2);
  assign _zz__13_7_inner_macOut_2 = (($signed(_zz__13_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_7_inner_activation;
    end else begin
      io_macOut = _13_7_inner_macOut;
    end
  end

  assign _zz__13_7_inner_macOut = ($signed(_zz__zz__13_7_inner_macOut) + $signed(_zz__zz__13_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_7_inner_activation <= 8'h00;
      _13_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_7_inner_activation <= io_addInput;
      end else begin
        _13_7_inner_macOut <= _zz__13_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_422 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_6_inner_macOut;
  wire       [15:0]   _zz__zz__13_6_inner_macOut_1;
  wire       [15:0]   _zz__13_6_inner_macOut_1;
  wire       [15:0]   _zz__13_6_inner_macOut_2;
  reg        [7:0]    _13_6_inner_activation;
  reg        [7:0]    _13_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_6_inner_macOut;

  assign _zz__zz__13_6_inner_macOut = ($signed(io_mulInput) * $signed(_13_6_inner_activation));
  assign _zz__zz__13_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_6_inner_macOut)) ? 16'h007f : _zz__13_6_inner_macOut_2);
  assign _zz__13_6_inner_macOut_2 = (($signed(_zz__13_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_6_inner_activation;
    end else begin
      io_macOut = _13_6_inner_macOut;
    end
  end

  assign _zz__13_6_inner_macOut = ($signed(_zz__zz__13_6_inner_macOut) + $signed(_zz__zz__13_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_6_inner_activation <= 8'h00;
      _13_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_6_inner_activation <= io_addInput;
      end else begin
        _13_6_inner_macOut <= _zz__13_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_421 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_5_inner_macOut;
  wire       [15:0]   _zz__zz__13_5_inner_macOut_1;
  wire       [15:0]   _zz__13_5_inner_macOut_1;
  wire       [15:0]   _zz__13_5_inner_macOut_2;
  reg        [7:0]    _13_5_inner_activation;
  reg        [7:0]    _13_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_5_inner_macOut;

  assign _zz__zz__13_5_inner_macOut = ($signed(io_mulInput) * $signed(_13_5_inner_activation));
  assign _zz__zz__13_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_5_inner_macOut)) ? 16'h007f : _zz__13_5_inner_macOut_2);
  assign _zz__13_5_inner_macOut_2 = (($signed(_zz__13_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_5_inner_activation;
    end else begin
      io_macOut = _13_5_inner_macOut;
    end
  end

  assign _zz__13_5_inner_macOut = ($signed(_zz__zz__13_5_inner_macOut) + $signed(_zz__zz__13_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_5_inner_activation <= 8'h00;
      _13_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_5_inner_activation <= io_addInput;
      end else begin
        _13_5_inner_macOut <= _zz__13_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_420 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_4_inner_macOut;
  wire       [15:0]   _zz__zz__13_4_inner_macOut_1;
  wire       [15:0]   _zz__13_4_inner_macOut_1;
  wire       [15:0]   _zz__13_4_inner_macOut_2;
  reg        [7:0]    _13_4_inner_activation;
  reg        [7:0]    _13_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_4_inner_macOut;

  assign _zz__zz__13_4_inner_macOut = ($signed(io_mulInput) * $signed(_13_4_inner_activation));
  assign _zz__zz__13_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_4_inner_macOut)) ? 16'h007f : _zz__13_4_inner_macOut_2);
  assign _zz__13_4_inner_macOut_2 = (($signed(_zz__13_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_4_inner_activation;
    end else begin
      io_macOut = _13_4_inner_macOut;
    end
  end

  assign _zz__13_4_inner_macOut = ($signed(_zz__zz__13_4_inner_macOut) + $signed(_zz__zz__13_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_4_inner_activation <= 8'h00;
      _13_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_4_inner_activation <= io_addInput;
      end else begin
        _13_4_inner_macOut <= _zz__13_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_419 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_3_inner_macOut;
  wire       [15:0]   _zz__zz__13_3_inner_macOut_1;
  wire       [15:0]   _zz__13_3_inner_macOut_1;
  wire       [15:0]   _zz__13_3_inner_macOut_2;
  reg        [7:0]    _13_3_inner_activation;
  reg        [7:0]    _13_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_3_inner_macOut;

  assign _zz__zz__13_3_inner_macOut = ($signed(io_mulInput) * $signed(_13_3_inner_activation));
  assign _zz__zz__13_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_3_inner_macOut)) ? 16'h007f : _zz__13_3_inner_macOut_2);
  assign _zz__13_3_inner_macOut_2 = (($signed(_zz__13_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_3_inner_activation;
    end else begin
      io_macOut = _13_3_inner_macOut;
    end
  end

  assign _zz__13_3_inner_macOut = ($signed(_zz__zz__13_3_inner_macOut) + $signed(_zz__zz__13_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_3_inner_activation <= 8'h00;
      _13_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_3_inner_activation <= io_addInput;
      end else begin
        _13_3_inner_macOut <= _zz__13_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_418 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_2_inner_macOut;
  wire       [15:0]   _zz__zz__13_2_inner_macOut_1;
  wire       [15:0]   _zz__13_2_inner_macOut_1;
  wire       [15:0]   _zz__13_2_inner_macOut_2;
  reg        [7:0]    _13_2_inner_activation;
  reg        [7:0]    _13_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_2_inner_macOut;

  assign _zz__zz__13_2_inner_macOut = ($signed(io_mulInput) * $signed(_13_2_inner_activation));
  assign _zz__zz__13_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_2_inner_macOut)) ? 16'h007f : _zz__13_2_inner_macOut_2);
  assign _zz__13_2_inner_macOut_2 = (($signed(_zz__13_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_2_inner_activation;
    end else begin
      io_macOut = _13_2_inner_macOut;
    end
  end

  assign _zz__13_2_inner_macOut = ($signed(_zz__zz__13_2_inner_macOut) + $signed(_zz__zz__13_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_2_inner_activation <= 8'h00;
      _13_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_2_inner_activation <= io_addInput;
      end else begin
        _13_2_inner_macOut <= _zz__13_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_417 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_1_inner_macOut;
  wire       [15:0]   _zz__zz__13_1_inner_macOut_1;
  wire       [15:0]   _zz__13_1_inner_macOut_1;
  wire       [15:0]   _zz__13_1_inner_macOut_2;
  reg        [7:0]    _13_1_inner_activation;
  reg        [7:0]    _13_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_1_inner_macOut;

  assign _zz__zz__13_1_inner_macOut = ($signed(io_mulInput) * $signed(_13_1_inner_activation));
  assign _zz__zz__13_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_1_inner_macOut)) ? 16'h007f : _zz__13_1_inner_macOut_2);
  assign _zz__13_1_inner_macOut_2 = (($signed(_zz__13_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_1_inner_activation;
    end else begin
      io_macOut = _13_1_inner_macOut;
    end
  end

  assign _zz__13_1_inner_macOut = ($signed(_zz__zz__13_1_inner_macOut) + $signed(_zz__zz__13_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_1_inner_activation <= 8'h00;
      _13_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_1_inner_activation <= io_addInput;
      end else begin
        _13_1_inner_macOut <= _zz__13_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_416 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__13_0_inner_macOut;
  wire       [15:0]   _zz__zz__13_0_inner_macOut_1;
  wire       [15:0]   _zz__13_0_inner_macOut_1;
  wire       [15:0]   _zz__13_0_inner_macOut_2;
  reg        [7:0]    _13_0_inner_activation;
  reg        [7:0]    _13_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__13_0_inner_macOut;

  assign _zz__zz__13_0_inner_macOut = ($signed(io_mulInput) * $signed(_13_0_inner_activation));
  assign _zz__zz__13_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__13_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__13_0_inner_macOut)) ? 16'h007f : _zz__13_0_inner_macOut_2);
  assign _zz__13_0_inner_macOut_2 = (($signed(_zz__13_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__13_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _13_0_inner_activation;
    end else begin
      io_macOut = _13_0_inner_macOut;
    end
  end

  assign _zz__13_0_inner_macOut = ($signed(_zz__zz__13_0_inner_macOut) + $signed(_zz__zz__13_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _13_0_inner_activation <= 8'h00;
      _13_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _13_0_inner_activation <= io_addInput;
      end else begin
        _13_0_inner_macOut <= _zz__13_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_415 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_31_inner_macOut;
  wire       [15:0]   _zz__zz__12_31_inner_macOut_1;
  wire       [15:0]   _zz__12_31_inner_macOut_1;
  wire       [15:0]   _zz__12_31_inner_macOut_2;
  reg        [7:0]    _12_31_inner_activation;
  reg        [7:0]    _12_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_31_inner_macOut;

  assign _zz__zz__12_31_inner_macOut = ($signed(io_mulInput) * $signed(_12_31_inner_activation));
  assign _zz__zz__12_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_31_inner_macOut)) ? 16'h007f : _zz__12_31_inner_macOut_2);
  assign _zz__12_31_inner_macOut_2 = (($signed(_zz__12_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_31_inner_activation;
    end else begin
      io_macOut = _12_31_inner_macOut;
    end
  end

  assign _zz__12_31_inner_macOut = ($signed(_zz__zz__12_31_inner_macOut) + $signed(_zz__zz__12_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_31_inner_activation <= 8'h00;
      _12_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_31_inner_activation <= io_addInput;
      end else begin
        _12_31_inner_macOut <= _zz__12_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_414 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_30_inner_macOut;
  wire       [15:0]   _zz__zz__12_30_inner_macOut_1;
  wire       [15:0]   _zz__12_30_inner_macOut_1;
  wire       [15:0]   _zz__12_30_inner_macOut_2;
  reg        [7:0]    _12_30_inner_activation;
  reg        [7:0]    _12_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_30_inner_macOut;

  assign _zz__zz__12_30_inner_macOut = ($signed(io_mulInput) * $signed(_12_30_inner_activation));
  assign _zz__zz__12_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_30_inner_macOut)) ? 16'h007f : _zz__12_30_inner_macOut_2);
  assign _zz__12_30_inner_macOut_2 = (($signed(_zz__12_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_30_inner_activation;
    end else begin
      io_macOut = _12_30_inner_macOut;
    end
  end

  assign _zz__12_30_inner_macOut = ($signed(_zz__zz__12_30_inner_macOut) + $signed(_zz__zz__12_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_30_inner_activation <= 8'h00;
      _12_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_30_inner_activation <= io_addInput;
      end else begin
        _12_30_inner_macOut <= _zz__12_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_413 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_29_inner_macOut;
  wire       [15:0]   _zz__zz__12_29_inner_macOut_1;
  wire       [15:0]   _zz__12_29_inner_macOut_1;
  wire       [15:0]   _zz__12_29_inner_macOut_2;
  reg        [7:0]    _12_29_inner_activation;
  reg        [7:0]    _12_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_29_inner_macOut;

  assign _zz__zz__12_29_inner_macOut = ($signed(io_mulInput) * $signed(_12_29_inner_activation));
  assign _zz__zz__12_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_29_inner_macOut)) ? 16'h007f : _zz__12_29_inner_macOut_2);
  assign _zz__12_29_inner_macOut_2 = (($signed(_zz__12_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_29_inner_activation;
    end else begin
      io_macOut = _12_29_inner_macOut;
    end
  end

  assign _zz__12_29_inner_macOut = ($signed(_zz__zz__12_29_inner_macOut) + $signed(_zz__zz__12_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_29_inner_activation <= 8'h00;
      _12_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_29_inner_activation <= io_addInput;
      end else begin
        _12_29_inner_macOut <= _zz__12_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_412 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_28_inner_macOut;
  wire       [15:0]   _zz__zz__12_28_inner_macOut_1;
  wire       [15:0]   _zz__12_28_inner_macOut_1;
  wire       [15:0]   _zz__12_28_inner_macOut_2;
  reg        [7:0]    _12_28_inner_activation;
  reg        [7:0]    _12_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_28_inner_macOut;

  assign _zz__zz__12_28_inner_macOut = ($signed(io_mulInput) * $signed(_12_28_inner_activation));
  assign _zz__zz__12_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_28_inner_macOut)) ? 16'h007f : _zz__12_28_inner_macOut_2);
  assign _zz__12_28_inner_macOut_2 = (($signed(_zz__12_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_28_inner_activation;
    end else begin
      io_macOut = _12_28_inner_macOut;
    end
  end

  assign _zz__12_28_inner_macOut = ($signed(_zz__zz__12_28_inner_macOut) + $signed(_zz__zz__12_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_28_inner_activation <= 8'h00;
      _12_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_28_inner_activation <= io_addInput;
      end else begin
        _12_28_inner_macOut <= _zz__12_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_411 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_27_inner_macOut;
  wire       [15:0]   _zz__zz__12_27_inner_macOut_1;
  wire       [15:0]   _zz__12_27_inner_macOut_1;
  wire       [15:0]   _zz__12_27_inner_macOut_2;
  reg        [7:0]    _12_27_inner_activation;
  reg        [7:0]    _12_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_27_inner_macOut;

  assign _zz__zz__12_27_inner_macOut = ($signed(io_mulInput) * $signed(_12_27_inner_activation));
  assign _zz__zz__12_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_27_inner_macOut)) ? 16'h007f : _zz__12_27_inner_macOut_2);
  assign _zz__12_27_inner_macOut_2 = (($signed(_zz__12_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_27_inner_activation;
    end else begin
      io_macOut = _12_27_inner_macOut;
    end
  end

  assign _zz__12_27_inner_macOut = ($signed(_zz__zz__12_27_inner_macOut) + $signed(_zz__zz__12_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_27_inner_activation <= 8'h00;
      _12_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_27_inner_activation <= io_addInput;
      end else begin
        _12_27_inner_macOut <= _zz__12_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_410 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_26_inner_macOut;
  wire       [15:0]   _zz__zz__12_26_inner_macOut_1;
  wire       [15:0]   _zz__12_26_inner_macOut_1;
  wire       [15:0]   _zz__12_26_inner_macOut_2;
  reg        [7:0]    _12_26_inner_activation;
  reg        [7:0]    _12_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_26_inner_macOut;

  assign _zz__zz__12_26_inner_macOut = ($signed(io_mulInput) * $signed(_12_26_inner_activation));
  assign _zz__zz__12_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_26_inner_macOut)) ? 16'h007f : _zz__12_26_inner_macOut_2);
  assign _zz__12_26_inner_macOut_2 = (($signed(_zz__12_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_26_inner_activation;
    end else begin
      io_macOut = _12_26_inner_macOut;
    end
  end

  assign _zz__12_26_inner_macOut = ($signed(_zz__zz__12_26_inner_macOut) + $signed(_zz__zz__12_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_26_inner_activation <= 8'h00;
      _12_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_26_inner_activation <= io_addInput;
      end else begin
        _12_26_inner_macOut <= _zz__12_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_409 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_25_inner_macOut;
  wire       [15:0]   _zz__zz__12_25_inner_macOut_1;
  wire       [15:0]   _zz__12_25_inner_macOut_1;
  wire       [15:0]   _zz__12_25_inner_macOut_2;
  reg        [7:0]    _12_25_inner_activation;
  reg        [7:0]    _12_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_25_inner_macOut;

  assign _zz__zz__12_25_inner_macOut = ($signed(io_mulInput) * $signed(_12_25_inner_activation));
  assign _zz__zz__12_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_25_inner_macOut)) ? 16'h007f : _zz__12_25_inner_macOut_2);
  assign _zz__12_25_inner_macOut_2 = (($signed(_zz__12_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_25_inner_activation;
    end else begin
      io_macOut = _12_25_inner_macOut;
    end
  end

  assign _zz__12_25_inner_macOut = ($signed(_zz__zz__12_25_inner_macOut) + $signed(_zz__zz__12_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_25_inner_activation <= 8'h00;
      _12_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_25_inner_activation <= io_addInput;
      end else begin
        _12_25_inner_macOut <= _zz__12_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_408 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_24_inner_macOut;
  wire       [15:0]   _zz__zz__12_24_inner_macOut_1;
  wire       [15:0]   _zz__12_24_inner_macOut_1;
  wire       [15:0]   _zz__12_24_inner_macOut_2;
  reg        [7:0]    _12_24_inner_activation;
  reg        [7:0]    _12_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_24_inner_macOut;

  assign _zz__zz__12_24_inner_macOut = ($signed(io_mulInput) * $signed(_12_24_inner_activation));
  assign _zz__zz__12_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_24_inner_macOut)) ? 16'h007f : _zz__12_24_inner_macOut_2);
  assign _zz__12_24_inner_macOut_2 = (($signed(_zz__12_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_24_inner_activation;
    end else begin
      io_macOut = _12_24_inner_macOut;
    end
  end

  assign _zz__12_24_inner_macOut = ($signed(_zz__zz__12_24_inner_macOut) + $signed(_zz__zz__12_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_24_inner_activation <= 8'h00;
      _12_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_24_inner_activation <= io_addInput;
      end else begin
        _12_24_inner_macOut <= _zz__12_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_407 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_23_inner_macOut;
  wire       [15:0]   _zz__zz__12_23_inner_macOut_1;
  wire       [15:0]   _zz__12_23_inner_macOut_1;
  wire       [15:0]   _zz__12_23_inner_macOut_2;
  reg        [7:0]    _12_23_inner_activation;
  reg        [7:0]    _12_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_23_inner_macOut;

  assign _zz__zz__12_23_inner_macOut = ($signed(io_mulInput) * $signed(_12_23_inner_activation));
  assign _zz__zz__12_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_23_inner_macOut)) ? 16'h007f : _zz__12_23_inner_macOut_2);
  assign _zz__12_23_inner_macOut_2 = (($signed(_zz__12_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_23_inner_activation;
    end else begin
      io_macOut = _12_23_inner_macOut;
    end
  end

  assign _zz__12_23_inner_macOut = ($signed(_zz__zz__12_23_inner_macOut) + $signed(_zz__zz__12_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_23_inner_activation <= 8'h00;
      _12_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_23_inner_activation <= io_addInput;
      end else begin
        _12_23_inner_macOut <= _zz__12_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_406 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_22_inner_macOut;
  wire       [15:0]   _zz__zz__12_22_inner_macOut_1;
  wire       [15:0]   _zz__12_22_inner_macOut_1;
  wire       [15:0]   _zz__12_22_inner_macOut_2;
  reg        [7:0]    _12_22_inner_activation;
  reg        [7:0]    _12_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_22_inner_macOut;

  assign _zz__zz__12_22_inner_macOut = ($signed(io_mulInput) * $signed(_12_22_inner_activation));
  assign _zz__zz__12_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_22_inner_macOut)) ? 16'h007f : _zz__12_22_inner_macOut_2);
  assign _zz__12_22_inner_macOut_2 = (($signed(_zz__12_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_22_inner_activation;
    end else begin
      io_macOut = _12_22_inner_macOut;
    end
  end

  assign _zz__12_22_inner_macOut = ($signed(_zz__zz__12_22_inner_macOut) + $signed(_zz__zz__12_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_22_inner_activation <= 8'h00;
      _12_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_22_inner_activation <= io_addInput;
      end else begin
        _12_22_inner_macOut <= _zz__12_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_405 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_21_inner_macOut;
  wire       [15:0]   _zz__zz__12_21_inner_macOut_1;
  wire       [15:0]   _zz__12_21_inner_macOut_1;
  wire       [15:0]   _zz__12_21_inner_macOut_2;
  reg        [7:0]    _12_21_inner_activation;
  reg        [7:0]    _12_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_21_inner_macOut;

  assign _zz__zz__12_21_inner_macOut = ($signed(io_mulInput) * $signed(_12_21_inner_activation));
  assign _zz__zz__12_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_21_inner_macOut)) ? 16'h007f : _zz__12_21_inner_macOut_2);
  assign _zz__12_21_inner_macOut_2 = (($signed(_zz__12_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_21_inner_activation;
    end else begin
      io_macOut = _12_21_inner_macOut;
    end
  end

  assign _zz__12_21_inner_macOut = ($signed(_zz__zz__12_21_inner_macOut) + $signed(_zz__zz__12_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_21_inner_activation <= 8'h00;
      _12_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_21_inner_activation <= io_addInput;
      end else begin
        _12_21_inner_macOut <= _zz__12_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_404 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_20_inner_macOut;
  wire       [15:0]   _zz__zz__12_20_inner_macOut_1;
  wire       [15:0]   _zz__12_20_inner_macOut_1;
  wire       [15:0]   _zz__12_20_inner_macOut_2;
  reg        [7:0]    _12_20_inner_activation;
  reg        [7:0]    _12_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_20_inner_macOut;

  assign _zz__zz__12_20_inner_macOut = ($signed(io_mulInput) * $signed(_12_20_inner_activation));
  assign _zz__zz__12_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_20_inner_macOut)) ? 16'h007f : _zz__12_20_inner_macOut_2);
  assign _zz__12_20_inner_macOut_2 = (($signed(_zz__12_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_20_inner_activation;
    end else begin
      io_macOut = _12_20_inner_macOut;
    end
  end

  assign _zz__12_20_inner_macOut = ($signed(_zz__zz__12_20_inner_macOut) + $signed(_zz__zz__12_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_20_inner_activation <= 8'h00;
      _12_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_20_inner_activation <= io_addInput;
      end else begin
        _12_20_inner_macOut <= _zz__12_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_403 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_19_inner_macOut;
  wire       [15:0]   _zz__zz__12_19_inner_macOut_1;
  wire       [15:0]   _zz__12_19_inner_macOut_1;
  wire       [15:0]   _zz__12_19_inner_macOut_2;
  reg        [7:0]    _12_19_inner_activation;
  reg        [7:0]    _12_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_19_inner_macOut;

  assign _zz__zz__12_19_inner_macOut = ($signed(io_mulInput) * $signed(_12_19_inner_activation));
  assign _zz__zz__12_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_19_inner_macOut)) ? 16'h007f : _zz__12_19_inner_macOut_2);
  assign _zz__12_19_inner_macOut_2 = (($signed(_zz__12_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_19_inner_activation;
    end else begin
      io_macOut = _12_19_inner_macOut;
    end
  end

  assign _zz__12_19_inner_macOut = ($signed(_zz__zz__12_19_inner_macOut) + $signed(_zz__zz__12_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_19_inner_activation <= 8'h00;
      _12_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_19_inner_activation <= io_addInput;
      end else begin
        _12_19_inner_macOut <= _zz__12_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_402 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_18_inner_macOut;
  wire       [15:0]   _zz__zz__12_18_inner_macOut_1;
  wire       [15:0]   _zz__12_18_inner_macOut_1;
  wire       [15:0]   _zz__12_18_inner_macOut_2;
  reg        [7:0]    _12_18_inner_activation;
  reg        [7:0]    _12_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_18_inner_macOut;

  assign _zz__zz__12_18_inner_macOut = ($signed(io_mulInput) * $signed(_12_18_inner_activation));
  assign _zz__zz__12_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_18_inner_macOut)) ? 16'h007f : _zz__12_18_inner_macOut_2);
  assign _zz__12_18_inner_macOut_2 = (($signed(_zz__12_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_18_inner_activation;
    end else begin
      io_macOut = _12_18_inner_macOut;
    end
  end

  assign _zz__12_18_inner_macOut = ($signed(_zz__zz__12_18_inner_macOut) + $signed(_zz__zz__12_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_18_inner_activation <= 8'h00;
      _12_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_18_inner_activation <= io_addInput;
      end else begin
        _12_18_inner_macOut <= _zz__12_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_401 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_17_inner_macOut;
  wire       [15:0]   _zz__zz__12_17_inner_macOut_1;
  wire       [15:0]   _zz__12_17_inner_macOut_1;
  wire       [15:0]   _zz__12_17_inner_macOut_2;
  reg        [7:0]    _12_17_inner_activation;
  reg        [7:0]    _12_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_17_inner_macOut;

  assign _zz__zz__12_17_inner_macOut = ($signed(io_mulInput) * $signed(_12_17_inner_activation));
  assign _zz__zz__12_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_17_inner_macOut)) ? 16'h007f : _zz__12_17_inner_macOut_2);
  assign _zz__12_17_inner_macOut_2 = (($signed(_zz__12_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_17_inner_activation;
    end else begin
      io_macOut = _12_17_inner_macOut;
    end
  end

  assign _zz__12_17_inner_macOut = ($signed(_zz__zz__12_17_inner_macOut) + $signed(_zz__zz__12_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_17_inner_activation <= 8'h00;
      _12_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_17_inner_activation <= io_addInput;
      end else begin
        _12_17_inner_macOut <= _zz__12_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_400 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_16_inner_macOut;
  wire       [15:0]   _zz__zz__12_16_inner_macOut_1;
  wire       [15:0]   _zz__12_16_inner_macOut_1;
  wire       [15:0]   _zz__12_16_inner_macOut_2;
  reg        [7:0]    _12_16_inner_activation;
  reg        [7:0]    _12_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_16_inner_macOut;

  assign _zz__zz__12_16_inner_macOut = ($signed(io_mulInput) * $signed(_12_16_inner_activation));
  assign _zz__zz__12_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_16_inner_macOut)) ? 16'h007f : _zz__12_16_inner_macOut_2);
  assign _zz__12_16_inner_macOut_2 = (($signed(_zz__12_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_16_inner_activation;
    end else begin
      io_macOut = _12_16_inner_macOut;
    end
  end

  assign _zz__12_16_inner_macOut = ($signed(_zz__zz__12_16_inner_macOut) + $signed(_zz__zz__12_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_16_inner_activation <= 8'h00;
      _12_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_16_inner_activation <= io_addInput;
      end else begin
        _12_16_inner_macOut <= _zz__12_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_399 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_15_inner_macOut;
  wire       [15:0]   _zz__zz__12_15_inner_macOut_1;
  wire       [15:0]   _zz__12_15_inner_macOut_1;
  wire       [15:0]   _zz__12_15_inner_macOut_2;
  reg        [7:0]    _12_15_inner_activation;
  reg        [7:0]    _12_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_15_inner_macOut;

  assign _zz__zz__12_15_inner_macOut = ($signed(io_mulInput) * $signed(_12_15_inner_activation));
  assign _zz__zz__12_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_15_inner_macOut)) ? 16'h007f : _zz__12_15_inner_macOut_2);
  assign _zz__12_15_inner_macOut_2 = (($signed(_zz__12_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_15_inner_activation;
    end else begin
      io_macOut = _12_15_inner_macOut;
    end
  end

  assign _zz__12_15_inner_macOut = ($signed(_zz__zz__12_15_inner_macOut) + $signed(_zz__zz__12_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_15_inner_activation <= 8'h00;
      _12_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_15_inner_activation <= io_addInput;
      end else begin
        _12_15_inner_macOut <= _zz__12_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_398 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_14_inner_macOut;
  wire       [15:0]   _zz__zz__12_14_inner_macOut_1;
  wire       [15:0]   _zz__12_14_inner_macOut_1;
  wire       [15:0]   _zz__12_14_inner_macOut_2;
  reg        [7:0]    _12_14_inner_activation;
  reg        [7:0]    _12_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_14_inner_macOut;

  assign _zz__zz__12_14_inner_macOut = ($signed(io_mulInput) * $signed(_12_14_inner_activation));
  assign _zz__zz__12_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_14_inner_macOut)) ? 16'h007f : _zz__12_14_inner_macOut_2);
  assign _zz__12_14_inner_macOut_2 = (($signed(_zz__12_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_14_inner_activation;
    end else begin
      io_macOut = _12_14_inner_macOut;
    end
  end

  assign _zz__12_14_inner_macOut = ($signed(_zz__zz__12_14_inner_macOut) + $signed(_zz__zz__12_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_14_inner_activation <= 8'h00;
      _12_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_14_inner_activation <= io_addInput;
      end else begin
        _12_14_inner_macOut <= _zz__12_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_397 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_13_inner_macOut;
  wire       [15:0]   _zz__zz__12_13_inner_macOut_1;
  wire       [15:0]   _zz__12_13_inner_macOut_1;
  wire       [15:0]   _zz__12_13_inner_macOut_2;
  reg        [7:0]    _12_13_inner_activation;
  reg        [7:0]    _12_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_13_inner_macOut;

  assign _zz__zz__12_13_inner_macOut = ($signed(io_mulInput) * $signed(_12_13_inner_activation));
  assign _zz__zz__12_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_13_inner_macOut)) ? 16'h007f : _zz__12_13_inner_macOut_2);
  assign _zz__12_13_inner_macOut_2 = (($signed(_zz__12_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_13_inner_activation;
    end else begin
      io_macOut = _12_13_inner_macOut;
    end
  end

  assign _zz__12_13_inner_macOut = ($signed(_zz__zz__12_13_inner_macOut) + $signed(_zz__zz__12_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_13_inner_activation <= 8'h00;
      _12_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_13_inner_activation <= io_addInput;
      end else begin
        _12_13_inner_macOut <= _zz__12_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_396 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_12_inner_macOut;
  wire       [15:0]   _zz__zz__12_12_inner_macOut_1;
  wire       [15:0]   _zz__12_12_inner_macOut_1;
  wire       [15:0]   _zz__12_12_inner_macOut_2;
  reg        [7:0]    _12_12_inner_activation;
  reg        [7:0]    _12_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_12_inner_macOut;

  assign _zz__zz__12_12_inner_macOut = ($signed(io_mulInput) * $signed(_12_12_inner_activation));
  assign _zz__zz__12_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_12_inner_macOut)) ? 16'h007f : _zz__12_12_inner_macOut_2);
  assign _zz__12_12_inner_macOut_2 = (($signed(_zz__12_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_12_inner_activation;
    end else begin
      io_macOut = _12_12_inner_macOut;
    end
  end

  assign _zz__12_12_inner_macOut = ($signed(_zz__zz__12_12_inner_macOut) + $signed(_zz__zz__12_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_12_inner_activation <= 8'h00;
      _12_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_12_inner_activation <= io_addInput;
      end else begin
        _12_12_inner_macOut <= _zz__12_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_395 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_11_inner_macOut;
  wire       [15:0]   _zz__zz__12_11_inner_macOut_1;
  wire       [15:0]   _zz__12_11_inner_macOut_1;
  wire       [15:0]   _zz__12_11_inner_macOut_2;
  reg        [7:0]    _12_11_inner_activation;
  reg        [7:0]    _12_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_11_inner_macOut;

  assign _zz__zz__12_11_inner_macOut = ($signed(io_mulInput) * $signed(_12_11_inner_activation));
  assign _zz__zz__12_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_11_inner_macOut)) ? 16'h007f : _zz__12_11_inner_macOut_2);
  assign _zz__12_11_inner_macOut_2 = (($signed(_zz__12_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_11_inner_activation;
    end else begin
      io_macOut = _12_11_inner_macOut;
    end
  end

  assign _zz__12_11_inner_macOut = ($signed(_zz__zz__12_11_inner_macOut) + $signed(_zz__zz__12_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_11_inner_activation <= 8'h00;
      _12_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_11_inner_activation <= io_addInput;
      end else begin
        _12_11_inner_macOut <= _zz__12_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_394 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_10_inner_macOut;
  wire       [15:0]   _zz__zz__12_10_inner_macOut_1;
  wire       [15:0]   _zz__12_10_inner_macOut_1;
  wire       [15:0]   _zz__12_10_inner_macOut_2;
  reg        [7:0]    _12_10_inner_activation;
  reg        [7:0]    _12_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_10_inner_macOut;

  assign _zz__zz__12_10_inner_macOut = ($signed(io_mulInput) * $signed(_12_10_inner_activation));
  assign _zz__zz__12_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_10_inner_macOut)) ? 16'h007f : _zz__12_10_inner_macOut_2);
  assign _zz__12_10_inner_macOut_2 = (($signed(_zz__12_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_10_inner_activation;
    end else begin
      io_macOut = _12_10_inner_macOut;
    end
  end

  assign _zz__12_10_inner_macOut = ($signed(_zz__zz__12_10_inner_macOut) + $signed(_zz__zz__12_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_10_inner_activation <= 8'h00;
      _12_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_10_inner_activation <= io_addInput;
      end else begin
        _12_10_inner_macOut <= _zz__12_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_393 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_9_inner_macOut;
  wire       [15:0]   _zz__zz__12_9_inner_macOut_1;
  wire       [15:0]   _zz__12_9_inner_macOut_1;
  wire       [15:0]   _zz__12_9_inner_macOut_2;
  reg        [7:0]    _12_9_inner_activation;
  reg        [7:0]    _12_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_9_inner_macOut;

  assign _zz__zz__12_9_inner_macOut = ($signed(io_mulInput) * $signed(_12_9_inner_activation));
  assign _zz__zz__12_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_9_inner_macOut)) ? 16'h007f : _zz__12_9_inner_macOut_2);
  assign _zz__12_9_inner_macOut_2 = (($signed(_zz__12_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_9_inner_activation;
    end else begin
      io_macOut = _12_9_inner_macOut;
    end
  end

  assign _zz__12_9_inner_macOut = ($signed(_zz__zz__12_9_inner_macOut) + $signed(_zz__zz__12_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_9_inner_activation <= 8'h00;
      _12_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_9_inner_activation <= io_addInput;
      end else begin
        _12_9_inner_macOut <= _zz__12_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_392 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_8_inner_macOut;
  wire       [15:0]   _zz__zz__12_8_inner_macOut_1;
  wire       [15:0]   _zz__12_8_inner_macOut_1;
  wire       [15:0]   _zz__12_8_inner_macOut_2;
  reg        [7:0]    _12_8_inner_activation;
  reg        [7:0]    _12_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_8_inner_macOut;

  assign _zz__zz__12_8_inner_macOut = ($signed(io_mulInput) * $signed(_12_8_inner_activation));
  assign _zz__zz__12_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_8_inner_macOut)) ? 16'h007f : _zz__12_8_inner_macOut_2);
  assign _zz__12_8_inner_macOut_2 = (($signed(_zz__12_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_8_inner_activation;
    end else begin
      io_macOut = _12_8_inner_macOut;
    end
  end

  assign _zz__12_8_inner_macOut = ($signed(_zz__zz__12_8_inner_macOut) + $signed(_zz__zz__12_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_8_inner_activation <= 8'h00;
      _12_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_8_inner_activation <= io_addInput;
      end else begin
        _12_8_inner_macOut <= _zz__12_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_391 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_7_inner_macOut;
  wire       [15:0]   _zz__zz__12_7_inner_macOut_1;
  wire       [15:0]   _zz__12_7_inner_macOut_1;
  wire       [15:0]   _zz__12_7_inner_macOut_2;
  reg        [7:0]    _12_7_inner_activation;
  reg        [7:0]    _12_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_7_inner_macOut;

  assign _zz__zz__12_7_inner_macOut = ($signed(io_mulInput) * $signed(_12_7_inner_activation));
  assign _zz__zz__12_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_7_inner_macOut)) ? 16'h007f : _zz__12_7_inner_macOut_2);
  assign _zz__12_7_inner_macOut_2 = (($signed(_zz__12_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_7_inner_activation;
    end else begin
      io_macOut = _12_7_inner_macOut;
    end
  end

  assign _zz__12_7_inner_macOut = ($signed(_zz__zz__12_7_inner_macOut) + $signed(_zz__zz__12_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_7_inner_activation <= 8'h00;
      _12_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_7_inner_activation <= io_addInput;
      end else begin
        _12_7_inner_macOut <= _zz__12_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_390 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_6_inner_macOut;
  wire       [15:0]   _zz__zz__12_6_inner_macOut_1;
  wire       [15:0]   _zz__12_6_inner_macOut_1;
  wire       [15:0]   _zz__12_6_inner_macOut_2;
  reg        [7:0]    _12_6_inner_activation;
  reg        [7:0]    _12_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_6_inner_macOut;

  assign _zz__zz__12_6_inner_macOut = ($signed(io_mulInput) * $signed(_12_6_inner_activation));
  assign _zz__zz__12_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_6_inner_macOut)) ? 16'h007f : _zz__12_6_inner_macOut_2);
  assign _zz__12_6_inner_macOut_2 = (($signed(_zz__12_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_6_inner_activation;
    end else begin
      io_macOut = _12_6_inner_macOut;
    end
  end

  assign _zz__12_6_inner_macOut = ($signed(_zz__zz__12_6_inner_macOut) + $signed(_zz__zz__12_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_6_inner_activation <= 8'h00;
      _12_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_6_inner_activation <= io_addInput;
      end else begin
        _12_6_inner_macOut <= _zz__12_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_389 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_5_inner_macOut;
  wire       [15:0]   _zz__zz__12_5_inner_macOut_1;
  wire       [15:0]   _zz__12_5_inner_macOut_1;
  wire       [15:0]   _zz__12_5_inner_macOut_2;
  reg        [7:0]    _12_5_inner_activation;
  reg        [7:0]    _12_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_5_inner_macOut;

  assign _zz__zz__12_5_inner_macOut = ($signed(io_mulInput) * $signed(_12_5_inner_activation));
  assign _zz__zz__12_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_5_inner_macOut)) ? 16'h007f : _zz__12_5_inner_macOut_2);
  assign _zz__12_5_inner_macOut_2 = (($signed(_zz__12_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_5_inner_activation;
    end else begin
      io_macOut = _12_5_inner_macOut;
    end
  end

  assign _zz__12_5_inner_macOut = ($signed(_zz__zz__12_5_inner_macOut) + $signed(_zz__zz__12_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_5_inner_activation <= 8'h00;
      _12_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_5_inner_activation <= io_addInput;
      end else begin
        _12_5_inner_macOut <= _zz__12_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_388 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_4_inner_macOut;
  wire       [15:0]   _zz__zz__12_4_inner_macOut_1;
  wire       [15:0]   _zz__12_4_inner_macOut_1;
  wire       [15:0]   _zz__12_4_inner_macOut_2;
  reg        [7:0]    _12_4_inner_activation;
  reg        [7:0]    _12_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_4_inner_macOut;

  assign _zz__zz__12_4_inner_macOut = ($signed(io_mulInput) * $signed(_12_4_inner_activation));
  assign _zz__zz__12_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_4_inner_macOut)) ? 16'h007f : _zz__12_4_inner_macOut_2);
  assign _zz__12_4_inner_macOut_2 = (($signed(_zz__12_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_4_inner_activation;
    end else begin
      io_macOut = _12_4_inner_macOut;
    end
  end

  assign _zz__12_4_inner_macOut = ($signed(_zz__zz__12_4_inner_macOut) + $signed(_zz__zz__12_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_4_inner_activation <= 8'h00;
      _12_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_4_inner_activation <= io_addInput;
      end else begin
        _12_4_inner_macOut <= _zz__12_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_387 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_3_inner_macOut;
  wire       [15:0]   _zz__zz__12_3_inner_macOut_1;
  wire       [15:0]   _zz__12_3_inner_macOut_1;
  wire       [15:0]   _zz__12_3_inner_macOut_2;
  reg        [7:0]    _12_3_inner_activation;
  reg        [7:0]    _12_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_3_inner_macOut;

  assign _zz__zz__12_3_inner_macOut = ($signed(io_mulInput) * $signed(_12_3_inner_activation));
  assign _zz__zz__12_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_3_inner_macOut)) ? 16'h007f : _zz__12_3_inner_macOut_2);
  assign _zz__12_3_inner_macOut_2 = (($signed(_zz__12_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_3_inner_activation;
    end else begin
      io_macOut = _12_3_inner_macOut;
    end
  end

  assign _zz__12_3_inner_macOut = ($signed(_zz__zz__12_3_inner_macOut) + $signed(_zz__zz__12_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_3_inner_activation <= 8'h00;
      _12_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_3_inner_activation <= io_addInput;
      end else begin
        _12_3_inner_macOut <= _zz__12_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_386 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_2_inner_macOut;
  wire       [15:0]   _zz__zz__12_2_inner_macOut_1;
  wire       [15:0]   _zz__12_2_inner_macOut_1;
  wire       [15:0]   _zz__12_2_inner_macOut_2;
  reg        [7:0]    _12_2_inner_activation;
  reg        [7:0]    _12_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_2_inner_macOut;

  assign _zz__zz__12_2_inner_macOut = ($signed(io_mulInput) * $signed(_12_2_inner_activation));
  assign _zz__zz__12_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_2_inner_macOut)) ? 16'h007f : _zz__12_2_inner_macOut_2);
  assign _zz__12_2_inner_macOut_2 = (($signed(_zz__12_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_2_inner_activation;
    end else begin
      io_macOut = _12_2_inner_macOut;
    end
  end

  assign _zz__12_2_inner_macOut = ($signed(_zz__zz__12_2_inner_macOut) + $signed(_zz__zz__12_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_2_inner_activation <= 8'h00;
      _12_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_2_inner_activation <= io_addInput;
      end else begin
        _12_2_inner_macOut <= _zz__12_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_385 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_1_inner_macOut;
  wire       [15:0]   _zz__zz__12_1_inner_macOut_1;
  wire       [15:0]   _zz__12_1_inner_macOut_1;
  wire       [15:0]   _zz__12_1_inner_macOut_2;
  reg        [7:0]    _12_1_inner_activation;
  reg        [7:0]    _12_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_1_inner_macOut;

  assign _zz__zz__12_1_inner_macOut = ($signed(io_mulInput) * $signed(_12_1_inner_activation));
  assign _zz__zz__12_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_1_inner_macOut)) ? 16'h007f : _zz__12_1_inner_macOut_2);
  assign _zz__12_1_inner_macOut_2 = (($signed(_zz__12_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_1_inner_activation;
    end else begin
      io_macOut = _12_1_inner_macOut;
    end
  end

  assign _zz__12_1_inner_macOut = ($signed(_zz__zz__12_1_inner_macOut) + $signed(_zz__zz__12_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_1_inner_activation <= 8'h00;
      _12_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_1_inner_activation <= io_addInput;
      end else begin
        _12_1_inner_macOut <= _zz__12_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_384 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__12_0_inner_macOut;
  wire       [15:0]   _zz__zz__12_0_inner_macOut_1;
  wire       [15:0]   _zz__12_0_inner_macOut_1;
  wire       [15:0]   _zz__12_0_inner_macOut_2;
  reg        [7:0]    _12_0_inner_activation;
  reg        [7:0]    _12_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__12_0_inner_macOut;

  assign _zz__zz__12_0_inner_macOut = ($signed(io_mulInput) * $signed(_12_0_inner_activation));
  assign _zz__zz__12_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__12_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__12_0_inner_macOut)) ? 16'h007f : _zz__12_0_inner_macOut_2);
  assign _zz__12_0_inner_macOut_2 = (($signed(_zz__12_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__12_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _12_0_inner_activation;
    end else begin
      io_macOut = _12_0_inner_macOut;
    end
  end

  assign _zz__12_0_inner_macOut = ($signed(_zz__zz__12_0_inner_macOut) + $signed(_zz__zz__12_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _12_0_inner_activation <= 8'h00;
      _12_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _12_0_inner_activation <= io_addInput;
      end else begin
        _12_0_inner_macOut <= _zz__12_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_383 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_31_inner_macOut;
  wire       [15:0]   _zz__zz__11_31_inner_macOut_1;
  wire       [15:0]   _zz__11_31_inner_macOut_1;
  wire       [15:0]   _zz__11_31_inner_macOut_2;
  reg        [7:0]    _11_31_inner_activation;
  reg        [7:0]    _11_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_31_inner_macOut;

  assign _zz__zz__11_31_inner_macOut = ($signed(io_mulInput) * $signed(_11_31_inner_activation));
  assign _zz__zz__11_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_31_inner_macOut)) ? 16'h007f : _zz__11_31_inner_macOut_2);
  assign _zz__11_31_inner_macOut_2 = (($signed(_zz__11_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_31_inner_activation;
    end else begin
      io_macOut = _11_31_inner_macOut;
    end
  end

  assign _zz__11_31_inner_macOut = ($signed(_zz__zz__11_31_inner_macOut) + $signed(_zz__zz__11_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_31_inner_activation <= 8'h00;
      _11_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_31_inner_activation <= io_addInput;
      end else begin
        _11_31_inner_macOut <= _zz__11_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_382 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_30_inner_macOut;
  wire       [15:0]   _zz__zz__11_30_inner_macOut_1;
  wire       [15:0]   _zz__11_30_inner_macOut_1;
  wire       [15:0]   _zz__11_30_inner_macOut_2;
  reg        [7:0]    _11_30_inner_activation;
  reg        [7:0]    _11_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_30_inner_macOut;

  assign _zz__zz__11_30_inner_macOut = ($signed(io_mulInput) * $signed(_11_30_inner_activation));
  assign _zz__zz__11_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_30_inner_macOut)) ? 16'h007f : _zz__11_30_inner_macOut_2);
  assign _zz__11_30_inner_macOut_2 = (($signed(_zz__11_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_30_inner_activation;
    end else begin
      io_macOut = _11_30_inner_macOut;
    end
  end

  assign _zz__11_30_inner_macOut = ($signed(_zz__zz__11_30_inner_macOut) + $signed(_zz__zz__11_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_30_inner_activation <= 8'h00;
      _11_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_30_inner_activation <= io_addInput;
      end else begin
        _11_30_inner_macOut <= _zz__11_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_381 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_29_inner_macOut;
  wire       [15:0]   _zz__zz__11_29_inner_macOut_1;
  wire       [15:0]   _zz__11_29_inner_macOut_1;
  wire       [15:0]   _zz__11_29_inner_macOut_2;
  reg        [7:0]    _11_29_inner_activation;
  reg        [7:0]    _11_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_29_inner_macOut;

  assign _zz__zz__11_29_inner_macOut = ($signed(io_mulInput) * $signed(_11_29_inner_activation));
  assign _zz__zz__11_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_29_inner_macOut)) ? 16'h007f : _zz__11_29_inner_macOut_2);
  assign _zz__11_29_inner_macOut_2 = (($signed(_zz__11_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_29_inner_activation;
    end else begin
      io_macOut = _11_29_inner_macOut;
    end
  end

  assign _zz__11_29_inner_macOut = ($signed(_zz__zz__11_29_inner_macOut) + $signed(_zz__zz__11_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_29_inner_activation <= 8'h00;
      _11_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_29_inner_activation <= io_addInput;
      end else begin
        _11_29_inner_macOut <= _zz__11_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_380 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_28_inner_macOut;
  wire       [15:0]   _zz__zz__11_28_inner_macOut_1;
  wire       [15:0]   _zz__11_28_inner_macOut_1;
  wire       [15:0]   _zz__11_28_inner_macOut_2;
  reg        [7:0]    _11_28_inner_activation;
  reg        [7:0]    _11_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_28_inner_macOut;

  assign _zz__zz__11_28_inner_macOut = ($signed(io_mulInput) * $signed(_11_28_inner_activation));
  assign _zz__zz__11_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_28_inner_macOut)) ? 16'h007f : _zz__11_28_inner_macOut_2);
  assign _zz__11_28_inner_macOut_2 = (($signed(_zz__11_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_28_inner_activation;
    end else begin
      io_macOut = _11_28_inner_macOut;
    end
  end

  assign _zz__11_28_inner_macOut = ($signed(_zz__zz__11_28_inner_macOut) + $signed(_zz__zz__11_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_28_inner_activation <= 8'h00;
      _11_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_28_inner_activation <= io_addInput;
      end else begin
        _11_28_inner_macOut <= _zz__11_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_379 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_27_inner_macOut;
  wire       [15:0]   _zz__zz__11_27_inner_macOut_1;
  wire       [15:0]   _zz__11_27_inner_macOut_1;
  wire       [15:0]   _zz__11_27_inner_macOut_2;
  reg        [7:0]    _11_27_inner_activation;
  reg        [7:0]    _11_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_27_inner_macOut;

  assign _zz__zz__11_27_inner_macOut = ($signed(io_mulInput) * $signed(_11_27_inner_activation));
  assign _zz__zz__11_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_27_inner_macOut)) ? 16'h007f : _zz__11_27_inner_macOut_2);
  assign _zz__11_27_inner_macOut_2 = (($signed(_zz__11_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_27_inner_activation;
    end else begin
      io_macOut = _11_27_inner_macOut;
    end
  end

  assign _zz__11_27_inner_macOut = ($signed(_zz__zz__11_27_inner_macOut) + $signed(_zz__zz__11_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_27_inner_activation <= 8'h00;
      _11_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_27_inner_activation <= io_addInput;
      end else begin
        _11_27_inner_macOut <= _zz__11_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_378 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_26_inner_macOut;
  wire       [15:0]   _zz__zz__11_26_inner_macOut_1;
  wire       [15:0]   _zz__11_26_inner_macOut_1;
  wire       [15:0]   _zz__11_26_inner_macOut_2;
  reg        [7:0]    _11_26_inner_activation;
  reg        [7:0]    _11_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_26_inner_macOut;

  assign _zz__zz__11_26_inner_macOut = ($signed(io_mulInput) * $signed(_11_26_inner_activation));
  assign _zz__zz__11_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_26_inner_macOut)) ? 16'h007f : _zz__11_26_inner_macOut_2);
  assign _zz__11_26_inner_macOut_2 = (($signed(_zz__11_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_26_inner_activation;
    end else begin
      io_macOut = _11_26_inner_macOut;
    end
  end

  assign _zz__11_26_inner_macOut = ($signed(_zz__zz__11_26_inner_macOut) + $signed(_zz__zz__11_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_26_inner_activation <= 8'h00;
      _11_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_26_inner_activation <= io_addInput;
      end else begin
        _11_26_inner_macOut <= _zz__11_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_377 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_25_inner_macOut;
  wire       [15:0]   _zz__zz__11_25_inner_macOut_1;
  wire       [15:0]   _zz__11_25_inner_macOut_1;
  wire       [15:0]   _zz__11_25_inner_macOut_2;
  reg        [7:0]    _11_25_inner_activation;
  reg        [7:0]    _11_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_25_inner_macOut;

  assign _zz__zz__11_25_inner_macOut = ($signed(io_mulInput) * $signed(_11_25_inner_activation));
  assign _zz__zz__11_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_25_inner_macOut)) ? 16'h007f : _zz__11_25_inner_macOut_2);
  assign _zz__11_25_inner_macOut_2 = (($signed(_zz__11_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_25_inner_activation;
    end else begin
      io_macOut = _11_25_inner_macOut;
    end
  end

  assign _zz__11_25_inner_macOut = ($signed(_zz__zz__11_25_inner_macOut) + $signed(_zz__zz__11_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_25_inner_activation <= 8'h00;
      _11_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_25_inner_activation <= io_addInput;
      end else begin
        _11_25_inner_macOut <= _zz__11_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_376 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_24_inner_macOut;
  wire       [15:0]   _zz__zz__11_24_inner_macOut_1;
  wire       [15:0]   _zz__11_24_inner_macOut_1;
  wire       [15:0]   _zz__11_24_inner_macOut_2;
  reg        [7:0]    _11_24_inner_activation;
  reg        [7:0]    _11_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_24_inner_macOut;

  assign _zz__zz__11_24_inner_macOut = ($signed(io_mulInput) * $signed(_11_24_inner_activation));
  assign _zz__zz__11_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_24_inner_macOut)) ? 16'h007f : _zz__11_24_inner_macOut_2);
  assign _zz__11_24_inner_macOut_2 = (($signed(_zz__11_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_24_inner_activation;
    end else begin
      io_macOut = _11_24_inner_macOut;
    end
  end

  assign _zz__11_24_inner_macOut = ($signed(_zz__zz__11_24_inner_macOut) + $signed(_zz__zz__11_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_24_inner_activation <= 8'h00;
      _11_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_24_inner_activation <= io_addInput;
      end else begin
        _11_24_inner_macOut <= _zz__11_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_375 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_23_inner_macOut;
  wire       [15:0]   _zz__zz__11_23_inner_macOut_1;
  wire       [15:0]   _zz__11_23_inner_macOut_1;
  wire       [15:0]   _zz__11_23_inner_macOut_2;
  reg        [7:0]    _11_23_inner_activation;
  reg        [7:0]    _11_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_23_inner_macOut;

  assign _zz__zz__11_23_inner_macOut = ($signed(io_mulInput) * $signed(_11_23_inner_activation));
  assign _zz__zz__11_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_23_inner_macOut)) ? 16'h007f : _zz__11_23_inner_macOut_2);
  assign _zz__11_23_inner_macOut_2 = (($signed(_zz__11_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_23_inner_activation;
    end else begin
      io_macOut = _11_23_inner_macOut;
    end
  end

  assign _zz__11_23_inner_macOut = ($signed(_zz__zz__11_23_inner_macOut) + $signed(_zz__zz__11_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_23_inner_activation <= 8'h00;
      _11_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_23_inner_activation <= io_addInput;
      end else begin
        _11_23_inner_macOut <= _zz__11_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_374 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_22_inner_macOut;
  wire       [15:0]   _zz__zz__11_22_inner_macOut_1;
  wire       [15:0]   _zz__11_22_inner_macOut_1;
  wire       [15:0]   _zz__11_22_inner_macOut_2;
  reg        [7:0]    _11_22_inner_activation;
  reg        [7:0]    _11_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_22_inner_macOut;

  assign _zz__zz__11_22_inner_macOut = ($signed(io_mulInput) * $signed(_11_22_inner_activation));
  assign _zz__zz__11_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_22_inner_macOut)) ? 16'h007f : _zz__11_22_inner_macOut_2);
  assign _zz__11_22_inner_macOut_2 = (($signed(_zz__11_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_22_inner_activation;
    end else begin
      io_macOut = _11_22_inner_macOut;
    end
  end

  assign _zz__11_22_inner_macOut = ($signed(_zz__zz__11_22_inner_macOut) + $signed(_zz__zz__11_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_22_inner_activation <= 8'h00;
      _11_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_22_inner_activation <= io_addInput;
      end else begin
        _11_22_inner_macOut <= _zz__11_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_373 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_21_inner_macOut;
  wire       [15:0]   _zz__zz__11_21_inner_macOut_1;
  wire       [15:0]   _zz__11_21_inner_macOut_1;
  wire       [15:0]   _zz__11_21_inner_macOut_2;
  reg        [7:0]    _11_21_inner_activation;
  reg        [7:0]    _11_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_21_inner_macOut;

  assign _zz__zz__11_21_inner_macOut = ($signed(io_mulInput) * $signed(_11_21_inner_activation));
  assign _zz__zz__11_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_21_inner_macOut)) ? 16'h007f : _zz__11_21_inner_macOut_2);
  assign _zz__11_21_inner_macOut_2 = (($signed(_zz__11_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_21_inner_activation;
    end else begin
      io_macOut = _11_21_inner_macOut;
    end
  end

  assign _zz__11_21_inner_macOut = ($signed(_zz__zz__11_21_inner_macOut) + $signed(_zz__zz__11_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_21_inner_activation <= 8'h00;
      _11_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_21_inner_activation <= io_addInput;
      end else begin
        _11_21_inner_macOut <= _zz__11_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_372 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_20_inner_macOut;
  wire       [15:0]   _zz__zz__11_20_inner_macOut_1;
  wire       [15:0]   _zz__11_20_inner_macOut_1;
  wire       [15:0]   _zz__11_20_inner_macOut_2;
  reg        [7:0]    _11_20_inner_activation;
  reg        [7:0]    _11_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_20_inner_macOut;

  assign _zz__zz__11_20_inner_macOut = ($signed(io_mulInput) * $signed(_11_20_inner_activation));
  assign _zz__zz__11_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_20_inner_macOut)) ? 16'h007f : _zz__11_20_inner_macOut_2);
  assign _zz__11_20_inner_macOut_2 = (($signed(_zz__11_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_20_inner_activation;
    end else begin
      io_macOut = _11_20_inner_macOut;
    end
  end

  assign _zz__11_20_inner_macOut = ($signed(_zz__zz__11_20_inner_macOut) + $signed(_zz__zz__11_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_20_inner_activation <= 8'h00;
      _11_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_20_inner_activation <= io_addInput;
      end else begin
        _11_20_inner_macOut <= _zz__11_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_371 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_19_inner_macOut;
  wire       [15:0]   _zz__zz__11_19_inner_macOut_1;
  wire       [15:0]   _zz__11_19_inner_macOut_1;
  wire       [15:0]   _zz__11_19_inner_macOut_2;
  reg        [7:0]    _11_19_inner_activation;
  reg        [7:0]    _11_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_19_inner_macOut;

  assign _zz__zz__11_19_inner_macOut = ($signed(io_mulInput) * $signed(_11_19_inner_activation));
  assign _zz__zz__11_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_19_inner_macOut)) ? 16'h007f : _zz__11_19_inner_macOut_2);
  assign _zz__11_19_inner_macOut_2 = (($signed(_zz__11_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_19_inner_activation;
    end else begin
      io_macOut = _11_19_inner_macOut;
    end
  end

  assign _zz__11_19_inner_macOut = ($signed(_zz__zz__11_19_inner_macOut) + $signed(_zz__zz__11_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_19_inner_activation <= 8'h00;
      _11_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_19_inner_activation <= io_addInput;
      end else begin
        _11_19_inner_macOut <= _zz__11_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_370 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_18_inner_macOut;
  wire       [15:0]   _zz__zz__11_18_inner_macOut_1;
  wire       [15:0]   _zz__11_18_inner_macOut_1;
  wire       [15:0]   _zz__11_18_inner_macOut_2;
  reg        [7:0]    _11_18_inner_activation;
  reg        [7:0]    _11_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_18_inner_macOut;

  assign _zz__zz__11_18_inner_macOut = ($signed(io_mulInput) * $signed(_11_18_inner_activation));
  assign _zz__zz__11_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_18_inner_macOut)) ? 16'h007f : _zz__11_18_inner_macOut_2);
  assign _zz__11_18_inner_macOut_2 = (($signed(_zz__11_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_18_inner_activation;
    end else begin
      io_macOut = _11_18_inner_macOut;
    end
  end

  assign _zz__11_18_inner_macOut = ($signed(_zz__zz__11_18_inner_macOut) + $signed(_zz__zz__11_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_18_inner_activation <= 8'h00;
      _11_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_18_inner_activation <= io_addInput;
      end else begin
        _11_18_inner_macOut <= _zz__11_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_369 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_17_inner_macOut;
  wire       [15:0]   _zz__zz__11_17_inner_macOut_1;
  wire       [15:0]   _zz__11_17_inner_macOut_1;
  wire       [15:0]   _zz__11_17_inner_macOut_2;
  reg        [7:0]    _11_17_inner_activation;
  reg        [7:0]    _11_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_17_inner_macOut;

  assign _zz__zz__11_17_inner_macOut = ($signed(io_mulInput) * $signed(_11_17_inner_activation));
  assign _zz__zz__11_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_17_inner_macOut)) ? 16'h007f : _zz__11_17_inner_macOut_2);
  assign _zz__11_17_inner_macOut_2 = (($signed(_zz__11_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_17_inner_activation;
    end else begin
      io_macOut = _11_17_inner_macOut;
    end
  end

  assign _zz__11_17_inner_macOut = ($signed(_zz__zz__11_17_inner_macOut) + $signed(_zz__zz__11_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_17_inner_activation <= 8'h00;
      _11_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_17_inner_activation <= io_addInput;
      end else begin
        _11_17_inner_macOut <= _zz__11_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_368 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_16_inner_macOut;
  wire       [15:0]   _zz__zz__11_16_inner_macOut_1;
  wire       [15:0]   _zz__11_16_inner_macOut_1;
  wire       [15:0]   _zz__11_16_inner_macOut_2;
  reg        [7:0]    _11_16_inner_activation;
  reg        [7:0]    _11_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_16_inner_macOut;

  assign _zz__zz__11_16_inner_macOut = ($signed(io_mulInput) * $signed(_11_16_inner_activation));
  assign _zz__zz__11_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_16_inner_macOut)) ? 16'h007f : _zz__11_16_inner_macOut_2);
  assign _zz__11_16_inner_macOut_2 = (($signed(_zz__11_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_16_inner_activation;
    end else begin
      io_macOut = _11_16_inner_macOut;
    end
  end

  assign _zz__11_16_inner_macOut = ($signed(_zz__zz__11_16_inner_macOut) + $signed(_zz__zz__11_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_16_inner_activation <= 8'h00;
      _11_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_16_inner_activation <= io_addInput;
      end else begin
        _11_16_inner_macOut <= _zz__11_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_367 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_15_inner_macOut;
  wire       [15:0]   _zz__zz__11_15_inner_macOut_1;
  wire       [15:0]   _zz__11_15_inner_macOut_1;
  wire       [15:0]   _zz__11_15_inner_macOut_2;
  reg        [7:0]    _11_15_inner_activation;
  reg        [7:0]    _11_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_15_inner_macOut;

  assign _zz__zz__11_15_inner_macOut = ($signed(io_mulInput) * $signed(_11_15_inner_activation));
  assign _zz__zz__11_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_15_inner_macOut)) ? 16'h007f : _zz__11_15_inner_macOut_2);
  assign _zz__11_15_inner_macOut_2 = (($signed(_zz__11_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_15_inner_activation;
    end else begin
      io_macOut = _11_15_inner_macOut;
    end
  end

  assign _zz__11_15_inner_macOut = ($signed(_zz__zz__11_15_inner_macOut) + $signed(_zz__zz__11_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_15_inner_activation <= 8'h00;
      _11_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_15_inner_activation <= io_addInput;
      end else begin
        _11_15_inner_macOut <= _zz__11_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_366 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_14_inner_macOut;
  wire       [15:0]   _zz__zz__11_14_inner_macOut_1;
  wire       [15:0]   _zz__11_14_inner_macOut_1;
  wire       [15:0]   _zz__11_14_inner_macOut_2;
  reg        [7:0]    _11_14_inner_activation;
  reg        [7:0]    _11_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_14_inner_macOut;

  assign _zz__zz__11_14_inner_macOut = ($signed(io_mulInput) * $signed(_11_14_inner_activation));
  assign _zz__zz__11_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_14_inner_macOut)) ? 16'h007f : _zz__11_14_inner_macOut_2);
  assign _zz__11_14_inner_macOut_2 = (($signed(_zz__11_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_14_inner_activation;
    end else begin
      io_macOut = _11_14_inner_macOut;
    end
  end

  assign _zz__11_14_inner_macOut = ($signed(_zz__zz__11_14_inner_macOut) + $signed(_zz__zz__11_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_14_inner_activation <= 8'h00;
      _11_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_14_inner_activation <= io_addInput;
      end else begin
        _11_14_inner_macOut <= _zz__11_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_365 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_13_inner_macOut;
  wire       [15:0]   _zz__zz__11_13_inner_macOut_1;
  wire       [15:0]   _zz__11_13_inner_macOut_1;
  wire       [15:0]   _zz__11_13_inner_macOut_2;
  reg        [7:0]    _11_13_inner_activation;
  reg        [7:0]    _11_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_13_inner_macOut;

  assign _zz__zz__11_13_inner_macOut = ($signed(io_mulInput) * $signed(_11_13_inner_activation));
  assign _zz__zz__11_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_13_inner_macOut)) ? 16'h007f : _zz__11_13_inner_macOut_2);
  assign _zz__11_13_inner_macOut_2 = (($signed(_zz__11_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_13_inner_activation;
    end else begin
      io_macOut = _11_13_inner_macOut;
    end
  end

  assign _zz__11_13_inner_macOut = ($signed(_zz__zz__11_13_inner_macOut) + $signed(_zz__zz__11_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_13_inner_activation <= 8'h00;
      _11_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_13_inner_activation <= io_addInput;
      end else begin
        _11_13_inner_macOut <= _zz__11_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_364 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_12_inner_macOut;
  wire       [15:0]   _zz__zz__11_12_inner_macOut_1;
  wire       [15:0]   _zz__11_12_inner_macOut_1;
  wire       [15:0]   _zz__11_12_inner_macOut_2;
  reg        [7:0]    _11_12_inner_activation;
  reg        [7:0]    _11_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_12_inner_macOut;

  assign _zz__zz__11_12_inner_macOut = ($signed(io_mulInput) * $signed(_11_12_inner_activation));
  assign _zz__zz__11_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_12_inner_macOut)) ? 16'h007f : _zz__11_12_inner_macOut_2);
  assign _zz__11_12_inner_macOut_2 = (($signed(_zz__11_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_12_inner_activation;
    end else begin
      io_macOut = _11_12_inner_macOut;
    end
  end

  assign _zz__11_12_inner_macOut = ($signed(_zz__zz__11_12_inner_macOut) + $signed(_zz__zz__11_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_12_inner_activation <= 8'h00;
      _11_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_12_inner_activation <= io_addInput;
      end else begin
        _11_12_inner_macOut <= _zz__11_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_363 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_11_inner_macOut;
  wire       [15:0]   _zz__zz__11_11_inner_macOut_1;
  wire       [15:0]   _zz__11_11_inner_macOut_1;
  wire       [15:0]   _zz__11_11_inner_macOut_2;
  reg        [7:0]    _11_11_inner_activation;
  reg        [7:0]    _11_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_11_inner_macOut;

  assign _zz__zz__11_11_inner_macOut = ($signed(io_mulInput) * $signed(_11_11_inner_activation));
  assign _zz__zz__11_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_11_inner_macOut)) ? 16'h007f : _zz__11_11_inner_macOut_2);
  assign _zz__11_11_inner_macOut_2 = (($signed(_zz__11_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_11_inner_activation;
    end else begin
      io_macOut = _11_11_inner_macOut;
    end
  end

  assign _zz__11_11_inner_macOut = ($signed(_zz__zz__11_11_inner_macOut) + $signed(_zz__zz__11_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_11_inner_activation <= 8'h00;
      _11_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_11_inner_activation <= io_addInput;
      end else begin
        _11_11_inner_macOut <= _zz__11_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_362 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_10_inner_macOut;
  wire       [15:0]   _zz__zz__11_10_inner_macOut_1;
  wire       [15:0]   _zz__11_10_inner_macOut_1;
  wire       [15:0]   _zz__11_10_inner_macOut_2;
  reg        [7:0]    _11_10_inner_activation;
  reg        [7:0]    _11_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_10_inner_macOut;

  assign _zz__zz__11_10_inner_macOut = ($signed(io_mulInput) * $signed(_11_10_inner_activation));
  assign _zz__zz__11_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_10_inner_macOut)) ? 16'h007f : _zz__11_10_inner_macOut_2);
  assign _zz__11_10_inner_macOut_2 = (($signed(_zz__11_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_10_inner_activation;
    end else begin
      io_macOut = _11_10_inner_macOut;
    end
  end

  assign _zz__11_10_inner_macOut = ($signed(_zz__zz__11_10_inner_macOut) + $signed(_zz__zz__11_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_10_inner_activation <= 8'h00;
      _11_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_10_inner_activation <= io_addInput;
      end else begin
        _11_10_inner_macOut <= _zz__11_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_361 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_9_inner_macOut;
  wire       [15:0]   _zz__zz__11_9_inner_macOut_1;
  wire       [15:0]   _zz__11_9_inner_macOut_1;
  wire       [15:0]   _zz__11_9_inner_macOut_2;
  reg        [7:0]    _11_9_inner_activation;
  reg        [7:0]    _11_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_9_inner_macOut;

  assign _zz__zz__11_9_inner_macOut = ($signed(io_mulInput) * $signed(_11_9_inner_activation));
  assign _zz__zz__11_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_9_inner_macOut)) ? 16'h007f : _zz__11_9_inner_macOut_2);
  assign _zz__11_9_inner_macOut_2 = (($signed(_zz__11_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_9_inner_activation;
    end else begin
      io_macOut = _11_9_inner_macOut;
    end
  end

  assign _zz__11_9_inner_macOut = ($signed(_zz__zz__11_9_inner_macOut) + $signed(_zz__zz__11_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_9_inner_activation <= 8'h00;
      _11_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_9_inner_activation <= io_addInput;
      end else begin
        _11_9_inner_macOut <= _zz__11_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_360 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_8_inner_macOut;
  wire       [15:0]   _zz__zz__11_8_inner_macOut_1;
  wire       [15:0]   _zz__11_8_inner_macOut_1;
  wire       [15:0]   _zz__11_8_inner_macOut_2;
  reg        [7:0]    _11_8_inner_activation;
  reg        [7:0]    _11_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_8_inner_macOut;

  assign _zz__zz__11_8_inner_macOut = ($signed(io_mulInput) * $signed(_11_8_inner_activation));
  assign _zz__zz__11_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_8_inner_macOut)) ? 16'h007f : _zz__11_8_inner_macOut_2);
  assign _zz__11_8_inner_macOut_2 = (($signed(_zz__11_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_8_inner_activation;
    end else begin
      io_macOut = _11_8_inner_macOut;
    end
  end

  assign _zz__11_8_inner_macOut = ($signed(_zz__zz__11_8_inner_macOut) + $signed(_zz__zz__11_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_8_inner_activation <= 8'h00;
      _11_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_8_inner_activation <= io_addInput;
      end else begin
        _11_8_inner_macOut <= _zz__11_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_359 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_7_inner_macOut;
  wire       [15:0]   _zz__zz__11_7_inner_macOut_1;
  wire       [15:0]   _zz__11_7_inner_macOut_1;
  wire       [15:0]   _zz__11_7_inner_macOut_2;
  reg        [7:0]    _11_7_inner_activation;
  reg        [7:0]    _11_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_7_inner_macOut;

  assign _zz__zz__11_7_inner_macOut = ($signed(io_mulInput) * $signed(_11_7_inner_activation));
  assign _zz__zz__11_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_7_inner_macOut)) ? 16'h007f : _zz__11_7_inner_macOut_2);
  assign _zz__11_7_inner_macOut_2 = (($signed(_zz__11_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_7_inner_activation;
    end else begin
      io_macOut = _11_7_inner_macOut;
    end
  end

  assign _zz__11_7_inner_macOut = ($signed(_zz__zz__11_7_inner_macOut) + $signed(_zz__zz__11_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_7_inner_activation <= 8'h00;
      _11_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_7_inner_activation <= io_addInput;
      end else begin
        _11_7_inner_macOut <= _zz__11_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_358 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_6_inner_macOut;
  wire       [15:0]   _zz__zz__11_6_inner_macOut_1;
  wire       [15:0]   _zz__11_6_inner_macOut_1;
  wire       [15:0]   _zz__11_6_inner_macOut_2;
  reg        [7:0]    _11_6_inner_activation;
  reg        [7:0]    _11_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_6_inner_macOut;

  assign _zz__zz__11_6_inner_macOut = ($signed(io_mulInput) * $signed(_11_6_inner_activation));
  assign _zz__zz__11_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_6_inner_macOut)) ? 16'h007f : _zz__11_6_inner_macOut_2);
  assign _zz__11_6_inner_macOut_2 = (($signed(_zz__11_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_6_inner_activation;
    end else begin
      io_macOut = _11_6_inner_macOut;
    end
  end

  assign _zz__11_6_inner_macOut = ($signed(_zz__zz__11_6_inner_macOut) + $signed(_zz__zz__11_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_6_inner_activation <= 8'h00;
      _11_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_6_inner_activation <= io_addInput;
      end else begin
        _11_6_inner_macOut <= _zz__11_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_357 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_5_inner_macOut;
  wire       [15:0]   _zz__zz__11_5_inner_macOut_1;
  wire       [15:0]   _zz__11_5_inner_macOut_1;
  wire       [15:0]   _zz__11_5_inner_macOut_2;
  reg        [7:0]    _11_5_inner_activation;
  reg        [7:0]    _11_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_5_inner_macOut;

  assign _zz__zz__11_5_inner_macOut = ($signed(io_mulInput) * $signed(_11_5_inner_activation));
  assign _zz__zz__11_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_5_inner_macOut)) ? 16'h007f : _zz__11_5_inner_macOut_2);
  assign _zz__11_5_inner_macOut_2 = (($signed(_zz__11_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_5_inner_activation;
    end else begin
      io_macOut = _11_5_inner_macOut;
    end
  end

  assign _zz__11_5_inner_macOut = ($signed(_zz__zz__11_5_inner_macOut) + $signed(_zz__zz__11_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_5_inner_activation <= 8'h00;
      _11_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_5_inner_activation <= io_addInput;
      end else begin
        _11_5_inner_macOut <= _zz__11_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_356 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_4_inner_macOut;
  wire       [15:0]   _zz__zz__11_4_inner_macOut_1;
  wire       [15:0]   _zz__11_4_inner_macOut_1;
  wire       [15:0]   _zz__11_4_inner_macOut_2;
  reg        [7:0]    _11_4_inner_activation;
  reg        [7:0]    _11_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_4_inner_macOut;

  assign _zz__zz__11_4_inner_macOut = ($signed(io_mulInput) * $signed(_11_4_inner_activation));
  assign _zz__zz__11_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_4_inner_macOut)) ? 16'h007f : _zz__11_4_inner_macOut_2);
  assign _zz__11_4_inner_macOut_2 = (($signed(_zz__11_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_4_inner_activation;
    end else begin
      io_macOut = _11_4_inner_macOut;
    end
  end

  assign _zz__11_4_inner_macOut = ($signed(_zz__zz__11_4_inner_macOut) + $signed(_zz__zz__11_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_4_inner_activation <= 8'h00;
      _11_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_4_inner_activation <= io_addInput;
      end else begin
        _11_4_inner_macOut <= _zz__11_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_355 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_3_inner_macOut;
  wire       [15:0]   _zz__zz__11_3_inner_macOut_1;
  wire       [15:0]   _zz__11_3_inner_macOut_1;
  wire       [15:0]   _zz__11_3_inner_macOut_2;
  reg        [7:0]    _11_3_inner_activation;
  reg        [7:0]    _11_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_3_inner_macOut;

  assign _zz__zz__11_3_inner_macOut = ($signed(io_mulInput) * $signed(_11_3_inner_activation));
  assign _zz__zz__11_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_3_inner_macOut)) ? 16'h007f : _zz__11_3_inner_macOut_2);
  assign _zz__11_3_inner_macOut_2 = (($signed(_zz__11_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_3_inner_activation;
    end else begin
      io_macOut = _11_3_inner_macOut;
    end
  end

  assign _zz__11_3_inner_macOut = ($signed(_zz__zz__11_3_inner_macOut) + $signed(_zz__zz__11_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_3_inner_activation <= 8'h00;
      _11_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_3_inner_activation <= io_addInput;
      end else begin
        _11_3_inner_macOut <= _zz__11_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_354 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_2_inner_macOut;
  wire       [15:0]   _zz__zz__11_2_inner_macOut_1;
  wire       [15:0]   _zz__11_2_inner_macOut_1;
  wire       [15:0]   _zz__11_2_inner_macOut_2;
  reg        [7:0]    _11_2_inner_activation;
  reg        [7:0]    _11_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_2_inner_macOut;

  assign _zz__zz__11_2_inner_macOut = ($signed(io_mulInput) * $signed(_11_2_inner_activation));
  assign _zz__zz__11_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_2_inner_macOut)) ? 16'h007f : _zz__11_2_inner_macOut_2);
  assign _zz__11_2_inner_macOut_2 = (($signed(_zz__11_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_2_inner_activation;
    end else begin
      io_macOut = _11_2_inner_macOut;
    end
  end

  assign _zz__11_2_inner_macOut = ($signed(_zz__zz__11_2_inner_macOut) + $signed(_zz__zz__11_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_2_inner_activation <= 8'h00;
      _11_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_2_inner_activation <= io_addInput;
      end else begin
        _11_2_inner_macOut <= _zz__11_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_353 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_1_inner_macOut;
  wire       [15:0]   _zz__zz__11_1_inner_macOut_1;
  wire       [15:0]   _zz__11_1_inner_macOut_1;
  wire       [15:0]   _zz__11_1_inner_macOut_2;
  reg        [7:0]    _11_1_inner_activation;
  reg        [7:0]    _11_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_1_inner_macOut;

  assign _zz__zz__11_1_inner_macOut = ($signed(io_mulInput) * $signed(_11_1_inner_activation));
  assign _zz__zz__11_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_1_inner_macOut)) ? 16'h007f : _zz__11_1_inner_macOut_2);
  assign _zz__11_1_inner_macOut_2 = (($signed(_zz__11_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_1_inner_activation;
    end else begin
      io_macOut = _11_1_inner_macOut;
    end
  end

  assign _zz__11_1_inner_macOut = ($signed(_zz__zz__11_1_inner_macOut) + $signed(_zz__zz__11_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_1_inner_activation <= 8'h00;
      _11_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_1_inner_activation <= io_addInput;
      end else begin
        _11_1_inner_macOut <= _zz__11_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_352 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__11_0_inner_macOut;
  wire       [15:0]   _zz__zz__11_0_inner_macOut_1;
  wire       [15:0]   _zz__11_0_inner_macOut_1;
  wire       [15:0]   _zz__11_0_inner_macOut_2;
  reg        [7:0]    _11_0_inner_activation;
  reg        [7:0]    _11_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__11_0_inner_macOut;

  assign _zz__zz__11_0_inner_macOut = ($signed(io_mulInput) * $signed(_11_0_inner_activation));
  assign _zz__zz__11_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__11_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__11_0_inner_macOut)) ? 16'h007f : _zz__11_0_inner_macOut_2);
  assign _zz__11_0_inner_macOut_2 = (($signed(_zz__11_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__11_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _11_0_inner_activation;
    end else begin
      io_macOut = _11_0_inner_macOut;
    end
  end

  assign _zz__11_0_inner_macOut = ($signed(_zz__zz__11_0_inner_macOut) + $signed(_zz__zz__11_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _11_0_inner_activation <= 8'h00;
      _11_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _11_0_inner_activation <= io_addInput;
      end else begin
        _11_0_inner_macOut <= _zz__11_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_351 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_31_inner_macOut;
  wire       [15:0]   _zz__zz__10_31_inner_macOut_1;
  wire       [15:0]   _zz__10_31_inner_macOut_1;
  wire       [15:0]   _zz__10_31_inner_macOut_2;
  reg        [7:0]    _10_31_inner_activation;
  reg        [7:0]    _10_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_31_inner_macOut;

  assign _zz__zz__10_31_inner_macOut = ($signed(io_mulInput) * $signed(_10_31_inner_activation));
  assign _zz__zz__10_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_31_inner_macOut)) ? 16'h007f : _zz__10_31_inner_macOut_2);
  assign _zz__10_31_inner_macOut_2 = (($signed(_zz__10_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_31_inner_activation;
    end else begin
      io_macOut = _10_31_inner_macOut;
    end
  end

  assign _zz__10_31_inner_macOut = ($signed(_zz__zz__10_31_inner_macOut) + $signed(_zz__zz__10_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_31_inner_activation <= 8'h00;
      _10_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_31_inner_activation <= io_addInput;
      end else begin
        _10_31_inner_macOut <= _zz__10_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_350 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_30_inner_macOut;
  wire       [15:0]   _zz__zz__10_30_inner_macOut_1;
  wire       [15:0]   _zz__10_30_inner_macOut_1;
  wire       [15:0]   _zz__10_30_inner_macOut_2;
  reg        [7:0]    _10_30_inner_activation;
  reg        [7:0]    _10_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_30_inner_macOut;

  assign _zz__zz__10_30_inner_macOut = ($signed(io_mulInput) * $signed(_10_30_inner_activation));
  assign _zz__zz__10_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_30_inner_macOut)) ? 16'h007f : _zz__10_30_inner_macOut_2);
  assign _zz__10_30_inner_macOut_2 = (($signed(_zz__10_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_30_inner_activation;
    end else begin
      io_macOut = _10_30_inner_macOut;
    end
  end

  assign _zz__10_30_inner_macOut = ($signed(_zz__zz__10_30_inner_macOut) + $signed(_zz__zz__10_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_30_inner_activation <= 8'h00;
      _10_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_30_inner_activation <= io_addInput;
      end else begin
        _10_30_inner_macOut <= _zz__10_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_349 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_29_inner_macOut;
  wire       [15:0]   _zz__zz__10_29_inner_macOut_1;
  wire       [15:0]   _zz__10_29_inner_macOut_1;
  wire       [15:0]   _zz__10_29_inner_macOut_2;
  reg        [7:0]    _10_29_inner_activation;
  reg        [7:0]    _10_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_29_inner_macOut;

  assign _zz__zz__10_29_inner_macOut = ($signed(io_mulInput) * $signed(_10_29_inner_activation));
  assign _zz__zz__10_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_29_inner_macOut)) ? 16'h007f : _zz__10_29_inner_macOut_2);
  assign _zz__10_29_inner_macOut_2 = (($signed(_zz__10_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_29_inner_activation;
    end else begin
      io_macOut = _10_29_inner_macOut;
    end
  end

  assign _zz__10_29_inner_macOut = ($signed(_zz__zz__10_29_inner_macOut) + $signed(_zz__zz__10_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_29_inner_activation <= 8'h00;
      _10_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_29_inner_activation <= io_addInput;
      end else begin
        _10_29_inner_macOut <= _zz__10_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_348 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_28_inner_macOut;
  wire       [15:0]   _zz__zz__10_28_inner_macOut_1;
  wire       [15:0]   _zz__10_28_inner_macOut_1;
  wire       [15:0]   _zz__10_28_inner_macOut_2;
  reg        [7:0]    _10_28_inner_activation;
  reg        [7:0]    _10_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_28_inner_macOut;

  assign _zz__zz__10_28_inner_macOut = ($signed(io_mulInput) * $signed(_10_28_inner_activation));
  assign _zz__zz__10_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_28_inner_macOut)) ? 16'h007f : _zz__10_28_inner_macOut_2);
  assign _zz__10_28_inner_macOut_2 = (($signed(_zz__10_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_28_inner_activation;
    end else begin
      io_macOut = _10_28_inner_macOut;
    end
  end

  assign _zz__10_28_inner_macOut = ($signed(_zz__zz__10_28_inner_macOut) + $signed(_zz__zz__10_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_28_inner_activation <= 8'h00;
      _10_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_28_inner_activation <= io_addInput;
      end else begin
        _10_28_inner_macOut <= _zz__10_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_347 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_27_inner_macOut;
  wire       [15:0]   _zz__zz__10_27_inner_macOut_1;
  wire       [15:0]   _zz__10_27_inner_macOut_1;
  wire       [15:0]   _zz__10_27_inner_macOut_2;
  reg        [7:0]    _10_27_inner_activation;
  reg        [7:0]    _10_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_27_inner_macOut;

  assign _zz__zz__10_27_inner_macOut = ($signed(io_mulInput) * $signed(_10_27_inner_activation));
  assign _zz__zz__10_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_27_inner_macOut)) ? 16'h007f : _zz__10_27_inner_macOut_2);
  assign _zz__10_27_inner_macOut_2 = (($signed(_zz__10_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_27_inner_activation;
    end else begin
      io_macOut = _10_27_inner_macOut;
    end
  end

  assign _zz__10_27_inner_macOut = ($signed(_zz__zz__10_27_inner_macOut) + $signed(_zz__zz__10_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_27_inner_activation <= 8'h00;
      _10_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_27_inner_activation <= io_addInput;
      end else begin
        _10_27_inner_macOut <= _zz__10_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_346 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_26_inner_macOut;
  wire       [15:0]   _zz__zz__10_26_inner_macOut_1;
  wire       [15:0]   _zz__10_26_inner_macOut_1;
  wire       [15:0]   _zz__10_26_inner_macOut_2;
  reg        [7:0]    _10_26_inner_activation;
  reg        [7:0]    _10_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_26_inner_macOut;

  assign _zz__zz__10_26_inner_macOut = ($signed(io_mulInput) * $signed(_10_26_inner_activation));
  assign _zz__zz__10_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_26_inner_macOut)) ? 16'h007f : _zz__10_26_inner_macOut_2);
  assign _zz__10_26_inner_macOut_2 = (($signed(_zz__10_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_26_inner_activation;
    end else begin
      io_macOut = _10_26_inner_macOut;
    end
  end

  assign _zz__10_26_inner_macOut = ($signed(_zz__zz__10_26_inner_macOut) + $signed(_zz__zz__10_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_26_inner_activation <= 8'h00;
      _10_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_26_inner_activation <= io_addInput;
      end else begin
        _10_26_inner_macOut <= _zz__10_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_345 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_25_inner_macOut;
  wire       [15:0]   _zz__zz__10_25_inner_macOut_1;
  wire       [15:0]   _zz__10_25_inner_macOut_1;
  wire       [15:0]   _zz__10_25_inner_macOut_2;
  reg        [7:0]    _10_25_inner_activation;
  reg        [7:0]    _10_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_25_inner_macOut;

  assign _zz__zz__10_25_inner_macOut = ($signed(io_mulInput) * $signed(_10_25_inner_activation));
  assign _zz__zz__10_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_25_inner_macOut)) ? 16'h007f : _zz__10_25_inner_macOut_2);
  assign _zz__10_25_inner_macOut_2 = (($signed(_zz__10_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_25_inner_activation;
    end else begin
      io_macOut = _10_25_inner_macOut;
    end
  end

  assign _zz__10_25_inner_macOut = ($signed(_zz__zz__10_25_inner_macOut) + $signed(_zz__zz__10_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_25_inner_activation <= 8'h00;
      _10_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_25_inner_activation <= io_addInput;
      end else begin
        _10_25_inner_macOut <= _zz__10_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_344 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_24_inner_macOut;
  wire       [15:0]   _zz__zz__10_24_inner_macOut_1;
  wire       [15:0]   _zz__10_24_inner_macOut_1;
  wire       [15:0]   _zz__10_24_inner_macOut_2;
  reg        [7:0]    _10_24_inner_activation;
  reg        [7:0]    _10_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_24_inner_macOut;

  assign _zz__zz__10_24_inner_macOut = ($signed(io_mulInput) * $signed(_10_24_inner_activation));
  assign _zz__zz__10_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_24_inner_macOut)) ? 16'h007f : _zz__10_24_inner_macOut_2);
  assign _zz__10_24_inner_macOut_2 = (($signed(_zz__10_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_24_inner_activation;
    end else begin
      io_macOut = _10_24_inner_macOut;
    end
  end

  assign _zz__10_24_inner_macOut = ($signed(_zz__zz__10_24_inner_macOut) + $signed(_zz__zz__10_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_24_inner_activation <= 8'h00;
      _10_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_24_inner_activation <= io_addInput;
      end else begin
        _10_24_inner_macOut <= _zz__10_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_343 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_23_inner_macOut;
  wire       [15:0]   _zz__zz__10_23_inner_macOut_1;
  wire       [15:0]   _zz__10_23_inner_macOut_1;
  wire       [15:0]   _zz__10_23_inner_macOut_2;
  reg        [7:0]    _10_23_inner_activation;
  reg        [7:0]    _10_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_23_inner_macOut;

  assign _zz__zz__10_23_inner_macOut = ($signed(io_mulInput) * $signed(_10_23_inner_activation));
  assign _zz__zz__10_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_23_inner_macOut)) ? 16'h007f : _zz__10_23_inner_macOut_2);
  assign _zz__10_23_inner_macOut_2 = (($signed(_zz__10_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_23_inner_activation;
    end else begin
      io_macOut = _10_23_inner_macOut;
    end
  end

  assign _zz__10_23_inner_macOut = ($signed(_zz__zz__10_23_inner_macOut) + $signed(_zz__zz__10_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_23_inner_activation <= 8'h00;
      _10_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_23_inner_activation <= io_addInput;
      end else begin
        _10_23_inner_macOut <= _zz__10_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_342 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_22_inner_macOut;
  wire       [15:0]   _zz__zz__10_22_inner_macOut_1;
  wire       [15:0]   _zz__10_22_inner_macOut_1;
  wire       [15:0]   _zz__10_22_inner_macOut_2;
  reg        [7:0]    _10_22_inner_activation;
  reg        [7:0]    _10_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_22_inner_macOut;

  assign _zz__zz__10_22_inner_macOut = ($signed(io_mulInput) * $signed(_10_22_inner_activation));
  assign _zz__zz__10_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_22_inner_macOut)) ? 16'h007f : _zz__10_22_inner_macOut_2);
  assign _zz__10_22_inner_macOut_2 = (($signed(_zz__10_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_22_inner_activation;
    end else begin
      io_macOut = _10_22_inner_macOut;
    end
  end

  assign _zz__10_22_inner_macOut = ($signed(_zz__zz__10_22_inner_macOut) + $signed(_zz__zz__10_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_22_inner_activation <= 8'h00;
      _10_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_22_inner_activation <= io_addInput;
      end else begin
        _10_22_inner_macOut <= _zz__10_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_341 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_21_inner_macOut;
  wire       [15:0]   _zz__zz__10_21_inner_macOut_1;
  wire       [15:0]   _zz__10_21_inner_macOut_1;
  wire       [15:0]   _zz__10_21_inner_macOut_2;
  reg        [7:0]    _10_21_inner_activation;
  reg        [7:0]    _10_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_21_inner_macOut;

  assign _zz__zz__10_21_inner_macOut = ($signed(io_mulInput) * $signed(_10_21_inner_activation));
  assign _zz__zz__10_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_21_inner_macOut)) ? 16'h007f : _zz__10_21_inner_macOut_2);
  assign _zz__10_21_inner_macOut_2 = (($signed(_zz__10_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_21_inner_activation;
    end else begin
      io_macOut = _10_21_inner_macOut;
    end
  end

  assign _zz__10_21_inner_macOut = ($signed(_zz__zz__10_21_inner_macOut) + $signed(_zz__zz__10_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_21_inner_activation <= 8'h00;
      _10_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_21_inner_activation <= io_addInput;
      end else begin
        _10_21_inner_macOut <= _zz__10_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_340 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_20_inner_macOut;
  wire       [15:0]   _zz__zz__10_20_inner_macOut_1;
  wire       [15:0]   _zz__10_20_inner_macOut_1;
  wire       [15:0]   _zz__10_20_inner_macOut_2;
  reg        [7:0]    _10_20_inner_activation;
  reg        [7:0]    _10_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_20_inner_macOut;

  assign _zz__zz__10_20_inner_macOut = ($signed(io_mulInput) * $signed(_10_20_inner_activation));
  assign _zz__zz__10_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_20_inner_macOut)) ? 16'h007f : _zz__10_20_inner_macOut_2);
  assign _zz__10_20_inner_macOut_2 = (($signed(_zz__10_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_20_inner_activation;
    end else begin
      io_macOut = _10_20_inner_macOut;
    end
  end

  assign _zz__10_20_inner_macOut = ($signed(_zz__zz__10_20_inner_macOut) + $signed(_zz__zz__10_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_20_inner_activation <= 8'h00;
      _10_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_20_inner_activation <= io_addInput;
      end else begin
        _10_20_inner_macOut <= _zz__10_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_339 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_19_inner_macOut;
  wire       [15:0]   _zz__zz__10_19_inner_macOut_1;
  wire       [15:0]   _zz__10_19_inner_macOut_1;
  wire       [15:0]   _zz__10_19_inner_macOut_2;
  reg        [7:0]    _10_19_inner_activation;
  reg        [7:0]    _10_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_19_inner_macOut;

  assign _zz__zz__10_19_inner_macOut = ($signed(io_mulInput) * $signed(_10_19_inner_activation));
  assign _zz__zz__10_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_19_inner_macOut)) ? 16'h007f : _zz__10_19_inner_macOut_2);
  assign _zz__10_19_inner_macOut_2 = (($signed(_zz__10_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_19_inner_activation;
    end else begin
      io_macOut = _10_19_inner_macOut;
    end
  end

  assign _zz__10_19_inner_macOut = ($signed(_zz__zz__10_19_inner_macOut) + $signed(_zz__zz__10_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_19_inner_activation <= 8'h00;
      _10_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_19_inner_activation <= io_addInput;
      end else begin
        _10_19_inner_macOut <= _zz__10_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_338 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_18_inner_macOut;
  wire       [15:0]   _zz__zz__10_18_inner_macOut_1;
  wire       [15:0]   _zz__10_18_inner_macOut_1;
  wire       [15:0]   _zz__10_18_inner_macOut_2;
  reg        [7:0]    _10_18_inner_activation;
  reg        [7:0]    _10_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_18_inner_macOut;

  assign _zz__zz__10_18_inner_macOut = ($signed(io_mulInput) * $signed(_10_18_inner_activation));
  assign _zz__zz__10_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_18_inner_macOut)) ? 16'h007f : _zz__10_18_inner_macOut_2);
  assign _zz__10_18_inner_macOut_2 = (($signed(_zz__10_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_18_inner_activation;
    end else begin
      io_macOut = _10_18_inner_macOut;
    end
  end

  assign _zz__10_18_inner_macOut = ($signed(_zz__zz__10_18_inner_macOut) + $signed(_zz__zz__10_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_18_inner_activation <= 8'h00;
      _10_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_18_inner_activation <= io_addInput;
      end else begin
        _10_18_inner_macOut <= _zz__10_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_337 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_17_inner_macOut;
  wire       [15:0]   _zz__zz__10_17_inner_macOut_1;
  wire       [15:0]   _zz__10_17_inner_macOut_1;
  wire       [15:0]   _zz__10_17_inner_macOut_2;
  reg        [7:0]    _10_17_inner_activation;
  reg        [7:0]    _10_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_17_inner_macOut;

  assign _zz__zz__10_17_inner_macOut = ($signed(io_mulInput) * $signed(_10_17_inner_activation));
  assign _zz__zz__10_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_17_inner_macOut)) ? 16'h007f : _zz__10_17_inner_macOut_2);
  assign _zz__10_17_inner_macOut_2 = (($signed(_zz__10_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_17_inner_activation;
    end else begin
      io_macOut = _10_17_inner_macOut;
    end
  end

  assign _zz__10_17_inner_macOut = ($signed(_zz__zz__10_17_inner_macOut) + $signed(_zz__zz__10_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_17_inner_activation <= 8'h00;
      _10_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_17_inner_activation <= io_addInput;
      end else begin
        _10_17_inner_macOut <= _zz__10_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_336 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_16_inner_macOut;
  wire       [15:0]   _zz__zz__10_16_inner_macOut_1;
  wire       [15:0]   _zz__10_16_inner_macOut_1;
  wire       [15:0]   _zz__10_16_inner_macOut_2;
  reg        [7:0]    _10_16_inner_activation;
  reg        [7:0]    _10_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_16_inner_macOut;

  assign _zz__zz__10_16_inner_macOut = ($signed(io_mulInput) * $signed(_10_16_inner_activation));
  assign _zz__zz__10_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_16_inner_macOut)) ? 16'h007f : _zz__10_16_inner_macOut_2);
  assign _zz__10_16_inner_macOut_2 = (($signed(_zz__10_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_16_inner_activation;
    end else begin
      io_macOut = _10_16_inner_macOut;
    end
  end

  assign _zz__10_16_inner_macOut = ($signed(_zz__zz__10_16_inner_macOut) + $signed(_zz__zz__10_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_16_inner_activation <= 8'h00;
      _10_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_16_inner_activation <= io_addInput;
      end else begin
        _10_16_inner_macOut <= _zz__10_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_335 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_15_inner_macOut;
  wire       [15:0]   _zz__zz__10_15_inner_macOut_1;
  wire       [15:0]   _zz__10_15_inner_macOut_1;
  wire       [15:0]   _zz__10_15_inner_macOut_2;
  reg        [7:0]    _10_15_inner_activation;
  reg        [7:0]    _10_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_15_inner_macOut;

  assign _zz__zz__10_15_inner_macOut = ($signed(io_mulInput) * $signed(_10_15_inner_activation));
  assign _zz__zz__10_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_15_inner_macOut)) ? 16'h007f : _zz__10_15_inner_macOut_2);
  assign _zz__10_15_inner_macOut_2 = (($signed(_zz__10_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_15_inner_activation;
    end else begin
      io_macOut = _10_15_inner_macOut;
    end
  end

  assign _zz__10_15_inner_macOut = ($signed(_zz__zz__10_15_inner_macOut) + $signed(_zz__zz__10_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_15_inner_activation <= 8'h00;
      _10_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_15_inner_activation <= io_addInput;
      end else begin
        _10_15_inner_macOut <= _zz__10_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_334 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_14_inner_macOut;
  wire       [15:0]   _zz__zz__10_14_inner_macOut_1;
  wire       [15:0]   _zz__10_14_inner_macOut_1;
  wire       [15:0]   _zz__10_14_inner_macOut_2;
  reg        [7:0]    _10_14_inner_activation;
  reg        [7:0]    _10_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_14_inner_macOut;

  assign _zz__zz__10_14_inner_macOut = ($signed(io_mulInput) * $signed(_10_14_inner_activation));
  assign _zz__zz__10_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_14_inner_macOut)) ? 16'h007f : _zz__10_14_inner_macOut_2);
  assign _zz__10_14_inner_macOut_2 = (($signed(_zz__10_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_14_inner_activation;
    end else begin
      io_macOut = _10_14_inner_macOut;
    end
  end

  assign _zz__10_14_inner_macOut = ($signed(_zz__zz__10_14_inner_macOut) + $signed(_zz__zz__10_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_14_inner_activation <= 8'h00;
      _10_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_14_inner_activation <= io_addInput;
      end else begin
        _10_14_inner_macOut <= _zz__10_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_333 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_13_inner_macOut;
  wire       [15:0]   _zz__zz__10_13_inner_macOut_1;
  wire       [15:0]   _zz__10_13_inner_macOut_1;
  wire       [15:0]   _zz__10_13_inner_macOut_2;
  reg        [7:0]    _10_13_inner_activation;
  reg        [7:0]    _10_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_13_inner_macOut;

  assign _zz__zz__10_13_inner_macOut = ($signed(io_mulInput) * $signed(_10_13_inner_activation));
  assign _zz__zz__10_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_13_inner_macOut)) ? 16'h007f : _zz__10_13_inner_macOut_2);
  assign _zz__10_13_inner_macOut_2 = (($signed(_zz__10_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_13_inner_activation;
    end else begin
      io_macOut = _10_13_inner_macOut;
    end
  end

  assign _zz__10_13_inner_macOut = ($signed(_zz__zz__10_13_inner_macOut) + $signed(_zz__zz__10_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_13_inner_activation <= 8'h00;
      _10_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_13_inner_activation <= io_addInput;
      end else begin
        _10_13_inner_macOut <= _zz__10_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_332 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_12_inner_macOut;
  wire       [15:0]   _zz__zz__10_12_inner_macOut_1;
  wire       [15:0]   _zz__10_12_inner_macOut_1;
  wire       [15:0]   _zz__10_12_inner_macOut_2;
  reg        [7:0]    _10_12_inner_activation;
  reg        [7:0]    _10_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_12_inner_macOut;

  assign _zz__zz__10_12_inner_macOut = ($signed(io_mulInput) * $signed(_10_12_inner_activation));
  assign _zz__zz__10_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_12_inner_macOut)) ? 16'h007f : _zz__10_12_inner_macOut_2);
  assign _zz__10_12_inner_macOut_2 = (($signed(_zz__10_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_12_inner_activation;
    end else begin
      io_macOut = _10_12_inner_macOut;
    end
  end

  assign _zz__10_12_inner_macOut = ($signed(_zz__zz__10_12_inner_macOut) + $signed(_zz__zz__10_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_12_inner_activation <= 8'h00;
      _10_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_12_inner_activation <= io_addInput;
      end else begin
        _10_12_inner_macOut <= _zz__10_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_331 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_11_inner_macOut;
  wire       [15:0]   _zz__zz__10_11_inner_macOut_1;
  wire       [15:0]   _zz__10_11_inner_macOut_1;
  wire       [15:0]   _zz__10_11_inner_macOut_2;
  reg        [7:0]    _10_11_inner_activation;
  reg        [7:0]    _10_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_11_inner_macOut;

  assign _zz__zz__10_11_inner_macOut = ($signed(io_mulInput) * $signed(_10_11_inner_activation));
  assign _zz__zz__10_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_11_inner_macOut)) ? 16'h007f : _zz__10_11_inner_macOut_2);
  assign _zz__10_11_inner_macOut_2 = (($signed(_zz__10_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_11_inner_activation;
    end else begin
      io_macOut = _10_11_inner_macOut;
    end
  end

  assign _zz__10_11_inner_macOut = ($signed(_zz__zz__10_11_inner_macOut) + $signed(_zz__zz__10_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_11_inner_activation <= 8'h00;
      _10_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_11_inner_activation <= io_addInput;
      end else begin
        _10_11_inner_macOut <= _zz__10_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_330 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_10_inner_macOut;
  wire       [15:0]   _zz__zz__10_10_inner_macOut_1;
  wire       [15:0]   _zz__10_10_inner_macOut_1;
  wire       [15:0]   _zz__10_10_inner_macOut_2;
  reg        [7:0]    _10_10_inner_activation;
  reg        [7:0]    _10_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_10_inner_macOut;

  assign _zz__zz__10_10_inner_macOut = ($signed(io_mulInput) * $signed(_10_10_inner_activation));
  assign _zz__zz__10_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_10_inner_macOut)) ? 16'h007f : _zz__10_10_inner_macOut_2);
  assign _zz__10_10_inner_macOut_2 = (($signed(_zz__10_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_10_inner_activation;
    end else begin
      io_macOut = _10_10_inner_macOut;
    end
  end

  assign _zz__10_10_inner_macOut = ($signed(_zz__zz__10_10_inner_macOut) + $signed(_zz__zz__10_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_10_inner_activation <= 8'h00;
      _10_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_10_inner_activation <= io_addInput;
      end else begin
        _10_10_inner_macOut <= _zz__10_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_329 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_9_inner_macOut;
  wire       [15:0]   _zz__zz__10_9_inner_macOut_1;
  wire       [15:0]   _zz__10_9_inner_macOut_1;
  wire       [15:0]   _zz__10_9_inner_macOut_2;
  reg        [7:0]    _10_9_inner_activation;
  reg        [7:0]    _10_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_9_inner_macOut;

  assign _zz__zz__10_9_inner_macOut = ($signed(io_mulInput) * $signed(_10_9_inner_activation));
  assign _zz__zz__10_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_9_inner_macOut)) ? 16'h007f : _zz__10_9_inner_macOut_2);
  assign _zz__10_9_inner_macOut_2 = (($signed(_zz__10_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_9_inner_activation;
    end else begin
      io_macOut = _10_9_inner_macOut;
    end
  end

  assign _zz__10_9_inner_macOut = ($signed(_zz__zz__10_9_inner_macOut) + $signed(_zz__zz__10_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_9_inner_activation <= 8'h00;
      _10_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_9_inner_activation <= io_addInput;
      end else begin
        _10_9_inner_macOut <= _zz__10_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_328 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_8_inner_macOut;
  wire       [15:0]   _zz__zz__10_8_inner_macOut_1;
  wire       [15:0]   _zz__10_8_inner_macOut_1;
  wire       [15:0]   _zz__10_8_inner_macOut_2;
  reg        [7:0]    _10_8_inner_activation;
  reg        [7:0]    _10_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_8_inner_macOut;

  assign _zz__zz__10_8_inner_macOut = ($signed(io_mulInput) * $signed(_10_8_inner_activation));
  assign _zz__zz__10_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_8_inner_macOut)) ? 16'h007f : _zz__10_8_inner_macOut_2);
  assign _zz__10_8_inner_macOut_2 = (($signed(_zz__10_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_8_inner_activation;
    end else begin
      io_macOut = _10_8_inner_macOut;
    end
  end

  assign _zz__10_8_inner_macOut = ($signed(_zz__zz__10_8_inner_macOut) + $signed(_zz__zz__10_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_8_inner_activation <= 8'h00;
      _10_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_8_inner_activation <= io_addInput;
      end else begin
        _10_8_inner_macOut <= _zz__10_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_327 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_7_inner_macOut;
  wire       [15:0]   _zz__zz__10_7_inner_macOut_1;
  wire       [15:0]   _zz__10_7_inner_macOut_1;
  wire       [15:0]   _zz__10_7_inner_macOut_2;
  reg        [7:0]    _10_7_inner_activation;
  reg        [7:0]    _10_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_7_inner_macOut;

  assign _zz__zz__10_7_inner_macOut = ($signed(io_mulInput) * $signed(_10_7_inner_activation));
  assign _zz__zz__10_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_7_inner_macOut)) ? 16'h007f : _zz__10_7_inner_macOut_2);
  assign _zz__10_7_inner_macOut_2 = (($signed(_zz__10_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_7_inner_activation;
    end else begin
      io_macOut = _10_7_inner_macOut;
    end
  end

  assign _zz__10_7_inner_macOut = ($signed(_zz__zz__10_7_inner_macOut) + $signed(_zz__zz__10_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_7_inner_activation <= 8'h00;
      _10_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_7_inner_activation <= io_addInput;
      end else begin
        _10_7_inner_macOut <= _zz__10_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_326 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_6_inner_macOut;
  wire       [15:0]   _zz__zz__10_6_inner_macOut_1;
  wire       [15:0]   _zz__10_6_inner_macOut_1;
  wire       [15:0]   _zz__10_6_inner_macOut_2;
  reg        [7:0]    _10_6_inner_activation;
  reg        [7:0]    _10_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_6_inner_macOut;

  assign _zz__zz__10_6_inner_macOut = ($signed(io_mulInput) * $signed(_10_6_inner_activation));
  assign _zz__zz__10_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_6_inner_macOut)) ? 16'h007f : _zz__10_6_inner_macOut_2);
  assign _zz__10_6_inner_macOut_2 = (($signed(_zz__10_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_6_inner_activation;
    end else begin
      io_macOut = _10_6_inner_macOut;
    end
  end

  assign _zz__10_6_inner_macOut = ($signed(_zz__zz__10_6_inner_macOut) + $signed(_zz__zz__10_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_6_inner_activation <= 8'h00;
      _10_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_6_inner_activation <= io_addInput;
      end else begin
        _10_6_inner_macOut <= _zz__10_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_325 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_5_inner_macOut;
  wire       [15:0]   _zz__zz__10_5_inner_macOut_1;
  wire       [15:0]   _zz__10_5_inner_macOut_1;
  wire       [15:0]   _zz__10_5_inner_macOut_2;
  reg        [7:0]    _10_5_inner_activation;
  reg        [7:0]    _10_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_5_inner_macOut;

  assign _zz__zz__10_5_inner_macOut = ($signed(io_mulInput) * $signed(_10_5_inner_activation));
  assign _zz__zz__10_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_5_inner_macOut)) ? 16'h007f : _zz__10_5_inner_macOut_2);
  assign _zz__10_5_inner_macOut_2 = (($signed(_zz__10_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_5_inner_activation;
    end else begin
      io_macOut = _10_5_inner_macOut;
    end
  end

  assign _zz__10_5_inner_macOut = ($signed(_zz__zz__10_5_inner_macOut) + $signed(_zz__zz__10_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_5_inner_activation <= 8'h00;
      _10_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_5_inner_activation <= io_addInput;
      end else begin
        _10_5_inner_macOut <= _zz__10_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_324 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_4_inner_macOut;
  wire       [15:0]   _zz__zz__10_4_inner_macOut_1;
  wire       [15:0]   _zz__10_4_inner_macOut_1;
  wire       [15:0]   _zz__10_4_inner_macOut_2;
  reg        [7:0]    _10_4_inner_activation;
  reg        [7:0]    _10_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_4_inner_macOut;

  assign _zz__zz__10_4_inner_macOut = ($signed(io_mulInput) * $signed(_10_4_inner_activation));
  assign _zz__zz__10_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_4_inner_macOut)) ? 16'h007f : _zz__10_4_inner_macOut_2);
  assign _zz__10_4_inner_macOut_2 = (($signed(_zz__10_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_4_inner_activation;
    end else begin
      io_macOut = _10_4_inner_macOut;
    end
  end

  assign _zz__10_4_inner_macOut = ($signed(_zz__zz__10_4_inner_macOut) + $signed(_zz__zz__10_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_4_inner_activation <= 8'h00;
      _10_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_4_inner_activation <= io_addInput;
      end else begin
        _10_4_inner_macOut <= _zz__10_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_323 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_3_inner_macOut;
  wire       [15:0]   _zz__zz__10_3_inner_macOut_1;
  wire       [15:0]   _zz__10_3_inner_macOut_1;
  wire       [15:0]   _zz__10_3_inner_macOut_2;
  reg        [7:0]    _10_3_inner_activation;
  reg        [7:0]    _10_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_3_inner_macOut;

  assign _zz__zz__10_3_inner_macOut = ($signed(io_mulInput) * $signed(_10_3_inner_activation));
  assign _zz__zz__10_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_3_inner_macOut)) ? 16'h007f : _zz__10_3_inner_macOut_2);
  assign _zz__10_3_inner_macOut_2 = (($signed(_zz__10_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_3_inner_activation;
    end else begin
      io_macOut = _10_3_inner_macOut;
    end
  end

  assign _zz__10_3_inner_macOut = ($signed(_zz__zz__10_3_inner_macOut) + $signed(_zz__zz__10_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_3_inner_activation <= 8'h00;
      _10_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_3_inner_activation <= io_addInput;
      end else begin
        _10_3_inner_macOut <= _zz__10_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_322 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_2_inner_macOut;
  wire       [15:0]   _zz__zz__10_2_inner_macOut_1;
  wire       [15:0]   _zz__10_2_inner_macOut_1;
  wire       [15:0]   _zz__10_2_inner_macOut_2;
  reg        [7:0]    _10_2_inner_activation;
  reg        [7:0]    _10_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_2_inner_macOut;

  assign _zz__zz__10_2_inner_macOut = ($signed(io_mulInput) * $signed(_10_2_inner_activation));
  assign _zz__zz__10_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_2_inner_macOut)) ? 16'h007f : _zz__10_2_inner_macOut_2);
  assign _zz__10_2_inner_macOut_2 = (($signed(_zz__10_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_2_inner_activation;
    end else begin
      io_macOut = _10_2_inner_macOut;
    end
  end

  assign _zz__10_2_inner_macOut = ($signed(_zz__zz__10_2_inner_macOut) + $signed(_zz__zz__10_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_2_inner_activation <= 8'h00;
      _10_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_2_inner_activation <= io_addInput;
      end else begin
        _10_2_inner_macOut <= _zz__10_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_321 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_1_inner_macOut;
  wire       [15:0]   _zz__zz__10_1_inner_macOut_1;
  wire       [15:0]   _zz__10_1_inner_macOut_1;
  wire       [15:0]   _zz__10_1_inner_macOut_2;
  reg        [7:0]    _10_1_inner_activation;
  reg        [7:0]    _10_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_1_inner_macOut;

  assign _zz__zz__10_1_inner_macOut = ($signed(io_mulInput) * $signed(_10_1_inner_activation));
  assign _zz__zz__10_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_1_inner_macOut)) ? 16'h007f : _zz__10_1_inner_macOut_2);
  assign _zz__10_1_inner_macOut_2 = (($signed(_zz__10_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_1_inner_activation;
    end else begin
      io_macOut = _10_1_inner_macOut;
    end
  end

  assign _zz__10_1_inner_macOut = ($signed(_zz__zz__10_1_inner_macOut) + $signed(_zz__zz__10_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_1_inner_activation <= 8'h00;
      _10_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_1_inner_activation <= io_addInput;
      end else begin
        _10_1_inner_macOut <= _zz__10_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_320 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__10_0_inner_macOut;
  wire       [15:0]   _zz__zz__10_0_inner_macOut_1;
  wire       [15:0]   _zz__10_0_inner_macOut_1;
  wire       [15:0]   _zz__10_0_inner_macOut_2;
  reg        [7:0]    _10_0_inner_activation;
  reg        [7:0]    _10_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__10_0_inner_macOut;

  assign _zz__zz__10_0_inner_macOut = ($signed(io_mulInput) * $signed(_10_0_inner_activation));
  assign _zz__zz__10_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__10_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__10_0_inner_macOut)) ? 16'h007f : _zz__10_0_inner_macOut_2);
  assign _zz__10_0_inner_macOut_2 = (($signed(_zz__10_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__10_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _10_0_inner_activation;
    end else begin
      io_macOut = _10_0_inner_macOut;
    end
  end

  assign _zz__10_0_inner_macOut = ($signed(_zz__zz__10_0_inner_macOut) + $signed(_zz__zz__10_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _10_0_inner_activation <= 8'h00;
      _10_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _10_0_inner_activation <= io_addInput;
      end else begin
        _10_0_inner_macOut <= _zz__10_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_319 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_31_inner_macOut;
  wire       [15:0]   _zz__zz__9_31_inner_macOut_1;
  wire       [15:0]   _zz__9_31_inner_macOut_1;
  wire       [15:0]   _zz__9_31_inner_macOut_2;
  reg        [7:0]    _9_31_inner_activation;
  reg        [7:0]    _9_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_31_inner_macOut;

  assign _zz__zz__9_31_inner_macOut = ($signed(io_mulInput) * $signed(_9_31_inner_activation));
  assign _zz__zz__9_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_31_inner_macOut)) ? 16'h007f : _zz__9_31_inner_macOut_2);
  assign _zz__9_31_inner_macOut_2 = (($signed(_zz__9_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_31_inner_activation;
    end else begin
      io_macOut = _9_31_inner_macOut;
    end
  end

  assign _zz__9_31_inner_macOut = ($signed(_zz__zz__9_31_inner_macOut) + $signed(_zz__zz__9_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_31_inner_activation <= 8'h00;
      _9_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_31_inner_activation <= io_addInput;
      end else begin
        _9_31_inner_macOut <= _zz__9_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_318 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_30_inner_macOut;
  wire       [15:0]   _zz__zz__9_30_inner_macOut_1;
  wire       [15:0]   _zz__9_30_inner_macOut_1;
  wire       [15:0]   _zz__9_30_inner_macOut_2;
  reg        [7:0]    _9_30_inner_activation;
  reg        [7:0]    _9_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_30_inner_macOut;

  assign _zz__zz__9_30_inner_macOut = ($signed(io_mulInput) * $signed(_9_30_inner_activation));
  assign _zz__zz__9_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_30_inner_macOut)) ? 16'h007f : _zz__9_30_inner_macOut_2);
  assign _zz__9_30_inner_macOut_2 = (($signed(_zz__9_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_30_inner_activation;
    end else begin
      io_macOut = _9_30_inner_macOut;
    end
  end

  assign _zz__9_30_inner_macOut = ($signed(_zz__zz__9_30_inner_macOut) + $signed(_zz__zz__9_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_30_inner_activation <= 8'h00;
      _9_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_30_inner_activation <= io_addInput;
      end else begin
        _9_30_inner_macOut <= _zz__9_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_317 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_29_inner_macOut;
  wire       [15:0]   _zz__zz__9_29_inner_macOut_1;
  wire       [15:0]   _zz__9_29_inner_macOut_1;
  wire       [15:0]   _zz__9_29_inner_macOut_2;
  reg        [7:0]    _9_29_inner_activation;
  reg        [7:0]    _9_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_29_inner_macOut;

  assign _zz__zz__9_29_inner_macOut = ($signed(io_mulInput) * $signed(_9_29_inner_activation));
  assign _zz__zz__9_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_29_inner_macOut)) ? 16'h007f : _zz__9_29_inner_macOut_2);
  assign _zz__9_29_inner_macOut_2 = (($signed(_zz__9_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_29_inner_activation;
    end else begin
      io_macOut = _9_29_inner_macOut;
    end
  end

  assign _zz__9_29_inner_macOut = ($signed(_zz__zz__9_29_inner_macOut) + $signed(_zz__zz__9_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_29_inner_activation <= 8'h00;
      _9_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_29_inner_activation <= io_addInput;
      end else begin
        _9_29_inner_macOut <= _zz__9_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_316 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_28_inner_macOut;
  wire       [15:0]   _zz__zz__9_28_inner_macOut_1;
  wire       [15:0]   _zz__9_28_inner_macOut_1;
  wire       [15:0]   _zz__9_28_inner_macOut_2;
  reg        [7:0]    _9_28_inner_activation;
  reg        [7:0]    _9_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_28_inner_macOut;

  assign _zz__zz__9_28_inner_macOut = ($signed(io_mulInput) * $signed(_9_28_inner_activation));
  assign _zz__zz__9_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_28_inner_macOut)) ? 16'h007f : _zz__9_28_inner_macOut_2);
  assign _zz__9_28_inner_macOut_2 = (($signed(_zz__9_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_28_inner_activation;
    end else begin
      io_macOut = _9_28_inner_macOut;
    end
  end

  assign _zz__9_28_inner_macOut = ($signed(_zz__zz__9_28_inner_macOut) + $signed(_zz__zz__9_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_28_inner_activation <= 8'h00;
      _9_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_28_inner_activation <= io_addInput;
      end else begin
        _9_28_inner_macOut <= _zz__9_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_315 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_27_inner_macOut;
  wire       [15:0]   _zz__zz__9_27_inner_macOut_1;
  wire       [15:0]   _zz__9_27_inner_macOut_1;
  wire       [15:0]   _zz__9_27_inner_macOut_2;
  reg        [7:0]    _9_27_inner_activation;
  reg        [7:0]    _9_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_27_inner_macOut;

  assign _zz__zz__9_27_inner_macOut = ($signed(io_mulInput) * $signed(_9_27_inner_activation));
  assign _zz__zz__9_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_27_inner_macOut)) ? 16'h007f : _zz__9_27_inner_macOut_2);
  assign _zz__9_27_inner_macOut_2 = (($signed(_zz__9_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_27_inner_activation;
    end else begin
      io_macOut = _9_27_inner_macOut;
    end
  end

  assign _zz__9_27_inner_macOut = ($signed(_zz__zz__9_27_inner_macOut) + $signed(_zz__zz__9_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_27_inner_activation <= 8'h00;
      _9_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_27_inner_activation <= io_addInput;
      end else begin
        _9_27_inner_macOut <= _zz__9_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_314 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_26_inner_macOut;
  wire       [15:0]   _zz__zz__9_26_inner_macOut_1;
  wire       [15:0]   _zz__9_26_inner_macOut_1;
  wire       [15:0]   _zz__9_26_inner_macOut_2;
  reg        [7:0]    _9_26_inner_activation;
  reg        [7:0]    _9_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_26_inner_macOut;

  assign _zz__zz__9_26_inner_macOut = ($signed(io_mulInput) * $signed(_9_26_inner_activation));
  assign _zz__zz__9_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_26_inner_macOut)) ? 16'h007f : _zz__9_26_inner_macOut_2);
  assign _zz__9_26_inner_macOut_2 = (($signed(_zz__9_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_26_inner_activation;
    end else begin
      io_macOut = _9_26_inner_macOut;
    end
  end

  assign _zz__9_26_inner_macOut = ($signed(_zz__zz__9_26_inner_macOut) + $signed(_zz__zz__9_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_26_inner_activation <= 8'h00;
      _9_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_26_inner_activation <= io_addInput;
      end else begin
        _9_26_inner_macOut <= _zz__9_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_313 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_25_inner_macOut;
  wire       [15:0]   _zz__zz__9_25_inner_macOut_1;
  wire       [15:0]   _zz__9_25_inner_macOut_1;
  wire       [15:0]   _zz__9_25_inner_macOut_2;
  reg        [7:0]    _9_25_inner_activation;
  reg        [7:0]    _9_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_25_inner_macOut;

  assign _zz__zz__9_25_inner_macOut = ($signed(io_mulInput) * $signed(_9_25_inner_activation));
  assign _zz__zz__9_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_25_inner_macOut)) ? 16'h007f : _zz__9_25_inner_macOut_2);
  assign _zz__9_25_inner_macOut_2 = (($signed(_zz__9_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_25_inner_activation;
    end else begin
      io_macOut = _9_25_inner_macOut;
    end
  end

  assign _zz__9_25_inner_macOut = ($signed(_zz__zz__9_25_inner_macOut) + $signed(_zz__zz__9_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_25_inner_activation <= 8'h00;
      _9_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_25_inner_activation <= io_addInput;
      end else begin
        _9_25_inner_macOut <= _zz__9_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_312 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_24_inner_macOut;
  wire       [15:0]   _zz__zz__9_24_inner_macOut_1;
  wire       [15:0]   _zz__9_24_inner_macOut_1;
  wire       [15:0]   _zz__9_24_inner_macOut_2;
  reg        [7:0]    _9_24_inner_activation;
  reg        [7:0]    _9_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_24_inner_macOut;

  assign _zz__zz__9_24_inner_macOut = ($signed(io_mulInput) * $signed(_9_24_inner_activation));
  assign _zz__zz__9_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_24_inner_macOut)) ? 16'h007f : _zz__9_24_inner_macOut_2);
  assign _zz__9_24_inner_macOut_2 = (($signed(_zz__9_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_24_inner_activation;
    end else begin
      io_macOut = _9_24_inner_macOut;
    end
  end

  assign _zz__9_24_inner_macOut = ($signed(_zz__zz__9_24_inner_macOut) + $signed(_zz__zz__9_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_24_inner_activation <= 8'h00;
      _9_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_24_inner_activation <= io_addInput;
      end else begin
        _9_24_inner_macOut <= _zz__9_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_311 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_23_inner_macOut;
  wire       [15:0]   _zz__zz__9_23_inner_macOut_1;
  wire       [15:0]   _zz__9_23_inner_macOut_1;
  wire       [15:0]   _zz__9_23_inner_macOut_2;
  reg        [7:0]    _9_23_inner_activation;
  reg        [7:0]    _9_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_23_inner_macOut;

  assign _zz__zz__9_23_inner_macOut = ($signed(io_mulInput) * $signed(_9_23_inner_activation));
  assign _zz__zz__9_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_23_inner_macOut)) ? 16'h007f : _zz__9_23_inner_macOut_2);
  assign _zz__9_23_inner_macOut_2 = (($signed(_zz__9_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_23_inner_activation;
    end else begin
      io_macOut = _9_23_inner_macOut;
    end
  end

  assign _zz__9_23_inner_macOut = ($signed(_zz__zz__9_23_inner_macOut) + $signed(_zz__zz__9_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_23_inner_activation <= 8'h00;
      _9_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_23_inner_activation <= io_addInput;
      end else begin
        _9_23_inner_macOut <= _zz__9_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_310 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_22_inner_macOut;
  wire       [15:0]   _zz__zz__9_22_inner_macOut_1;
  wire       [15:0]   _zz__9_22_inner_macOut_1;
  wire       [15:0]   _zz__9_22_inner_macOut_2;
  reg        [7:0]    _9_22_inner_activation;
  reg        [7:0]    _9_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_22_inner_macOut;

  assign _zz__zz__9_22_inner_macOut = ($signed(io_mulInput) * $signed(_9_22_inner_activation));
  assign _zz__zz__9_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_22_inner_macOut)) ? 16'h007f : _zz__9_22_inner_macOut_2);
  assign _zz__9_22_inner_macOut_2 = (($signed(_zz__9_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_22_inner_activation;
    end else begin
      io_macOut = _9_22_inner_macOut;
    end
  end

  assign _zz__9_22_inner_macOut = ($signed(_zz__zz__9_22_inner_macOut) + $signed(_zz__zz__9_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_22_inner_activation <= 8'h00;
      _9_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_22_inner_activation <= io_addInput;
      end else begin
        _9_22_inner_macOut <= _zz__9_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_309 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_21_inner_macOut;
  wire       [15:0]   _zz__zz__9_21_inner_macOut_1;
  wire       [15:0]   _zz__9_21_inner_macOut_1;
  wire       [15:0]   _zz__9_21_inner_macOut_2;
  reg        [7:0]    _9_21_inner_activation;
  reg        [7:0]    _9_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_21_inner_macOut;

  assign _zz__zz__9_21_inner_macOut = ($signed(io_mulInput) * $signed(_9_21_inner_activation));
  assign _zz__zz__9_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_21_inner_macOut)) ? 16'h007f : _zz__9_21_inner_macOut_2);
  assign _zz__9_21_inner_macOut_2 = (($signed(_zz__9_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_21_inner_activation;
    end else begin
      io_macOut = _9_21_inner_macOut;
    end
  end

  assign _zz__9_21_inner_macOut = ($signed(_zz__zz__9_21_inner_macOut) + $signed(_zz__zz__9_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_21_inner_activation <= 8'h00;
      _9_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_21_inner_activation <= io_addInput;
      end else begin
        _9_21_inner_macOut <= _zz__9_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_308 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_20_inner_macOut;
  wire       [15:0]   _zz__zz__9_20_inner_macOut_1;
  wire       [15:0]   _zz__9_20_inner_macOut_1;
  wire       [15:0]   _zz__9_20_inner_macOut_2;
  reg        [7:0]    _9_20_inner_activation;
  reg        [7:0]    _9_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_20_inner_macOut;

  assign _zz__zz__9_20_inner_macOut = ($signed(io_mulInput) * $signed(_9_20_inner_activation));
  assign _zz__zz__9_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_20_inner_macOut)) ? 16'h007f : _zz__9_20_inner_macOut_2);
  assign _zz__9_20_inner_macOut_2 = (($signed(_zz__9_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_20_inner_activation;
    end else begin
      io_macOut = _9_20_inner_macOut;
    end
  end

  assign _zz__9_20_inner_macOut = ($signed(_zz__zz__9_20_inner_macOut) + $signed(_zz__zz__9_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_20_inner_activation <= 8'h00;
      _9_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_20_inner_activation <= io_addInput;
      end else begin
        _9_20_inner_macOut <= _zz__9_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_307 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_19_inner_macOut;
  wire       [15:0]   _zz__zz__9_19_inner_macOut_1;
  wire       [15:0]   _zz__9_19_inner_macOut_1;
  wire       [15:0]   _zz__9_19_inner_macOut_2;
  reg        [7:0]    _9_19_inner_activation;
  reg        [7:0]    _9_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_19_inner_macOut;

  assign _zz__zz__9_19_inner_macOut = ($signed(io_mulInput) * $signed(_9_19_inner_activation));
  assign _zz__zz__9_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_19_inner_macOut)) ? 16'h007f : _zz__9_19_inner_macOut_2);
  assign _zz__9_19_inner_macOut_2 = (($signed(_zz__9_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_19_inner_activation;
    end else begin
      io_macOut = _9_19_inner_macOut;
    end
  end

  assign _zz__9_19_inner_macOut = ($signed(_zz__zz__9_19_inner_macOut) + $signed(_zz__zz__9_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_19_inner_activation <= 8'h00;
      _9_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_19_inner_activation <= io_addInput;
      end else begin
        _9_19_inner_macOut <= _zz__9_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_306 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_18_inner_macOut;
  wire       [15:0]   _zz__zz__9_18_inner_macOut_1;
  wire       [15:0]   _zz__9_18_inner_macOut_1;
  wire       [15:0]   _zz__9_18_inner_macOut_2;
  reg        [7:0]    _9_18_inner_activation;
  reg        [7:0]    _9_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_18_inner_macOut;

  assign _zz__zz__9_18_inner_macOut = ($signed(io_mulInput) * $signed(_9_18_inner_activation));
  assign _zz__zz__9_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_18_inner_macOut)) ? 16'h007f : _zz__9_18_inner_macOut_2);
  assign _zz__9_18_inner_macOut_2 = (($signed(_zz__9_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_18_inner_activation;
    end else begin
      io_macOut = _9_18_inner_macOut;
    end
  end

  assign _zz__9_18_inner_macOut = ($signed(_zz__zz__9_18_inner_macOut) + $signed(_zz__zz__9_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_18_inner_activation <= 8'h00;
      _9_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_18_inner_activation <= io_addInput;
      end else begin
        _9_18_inner_macOut <= _zz__9_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_305 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_17_inner_macOut;
  wire       [15:0]   _zz__zz__9_17_inner_macOut_1;
  wire       [15:0]   _zz__9_17_inner_macOut_1;
  wire       [15:0]   _zz__9_17_inner_macOut_2;
  reg        [7:0]    _9_17_inner_activation;
  reg        [7:0]    _9_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_17_inner_macOut;

  assign _zz__zz__9_17_inner_macOut = ($signed(io_mulInput) * $signed(_9_17_inner_activation));
  assign _zz__zz__9_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_17_inner_macOut)) ? 16'h007f : _zz__9_17_inner_macOut_2);
  assign _zz__9_17_inner_macOut_2 = (($signed(_zz__9_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_17_inner_activation;
    end else begin
      io_macOut = _9_17_inner_macOut;
    end
  end

  assign _zz__9_17_inner_macOut = ($signed(_zz__zz__9_17_inner_macOut) + $signed(_zz__zz__9_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_17_inner_activation <= 8'h00;
      _9_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_17_inner_activation <= io_addInput;
      end else begin
        _9_17_inner_macOut <= _zz__9_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_304 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_16_inner_macOut;
  wire       [15:0]   _zz__zz__9_16_inner_macOut_1;
  wire       [15:0]   _zz__9_16_inner_macOut_1;
  wire       [15:0]   _zz__9_16_inner_macOut_2;
  reg        [7:0]    _9_16_inner_activation;
  reg        [7:0]    _9_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_16_inner_macOut;

  assign _zz__zz__9_16_inner_macOut = ($signed(io_mulInput) * $signed(_9_16_inner_activation));
  assign _zz__zz__9_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_16_inner_macOut)) ? 16'h007f : _zz__9_16_inner_macOut_2);
  assign _zz__9_16_inner_macOut_2 = (($signed(_zz__9_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_16_inner_activation;
    end else begin
      io_macOut = _9_16_inner_macOut;
    end
  end

  assign _zz__9_16_inner_macOut = ($signed(_zz__zz__9_16_inner_macOut) + $signed(_zz__zz__9_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_16_inner_activation <= 8'h00;
      _9_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_16_inner_activation <= io_addInput;
      end else begin
        _9_16_inner_macOut <= _zz__9_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_303 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_15_inner_macOut;
  wire       [15:0]   _zz__zz__9_15_inner_macOut_1;
  wire       [15:0]   _zz__9_15_inner_macOut_1;
  wire       [15:0]   _zz__9_15_inner_macOut_2;
  reg        [7:0]    _9_15_inner_activation;
  reg        [7:0]    _9_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_15_inner_macOut;

  assign _zz__zz__9_15_inner_macOut = ($signed(io_mulInput) * $signed(_9_15_inner_activation));
  assign _zz__zz__9_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_15_inner_macOut)) ? 16'h007f : _zz__9_15_inner_macOut_2);
  assign _zz__9_15_inner_macOut_2 = (($signed(_zz__9_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_15_inner_activation;
    end else begin
      io_macOut = _9_15_inner_macOut;
    end
  end

  assign _zz__9_15_inner_macOut = ($signed(_zz__zz__9_15_inner_macOut) + $signed(_zz__zz__9_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_15_inner_activation <= 8'h00;
      _9_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_15_inner_activation <= io_addInput;
      end else begin
        _9_15_inner_macOut <= _zz__9_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_302 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_14_inner_macOut;
  wire       [15:0]   _zz__zz__9_14_inner_macOut_1;
  wire       [15:0]   _zz__9_14_inner_macOut_1;
  wire       [15:0]   _zz__9_14_inner_macOut_2;
  reg        [7:0]    _9_14_inner_activation;
  reg        [7:0]    _9_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_14_inner_macOut;

  assign _zz__zz__9_14_inner_macOut = ($signed(io_mulInput) * $signed(_9_14_inner_activation));
  assign _zz__zz__9_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_14_inner_macOut)) ? 16'h007f : _zz__9_14_inner_macOut_2);
  assign _zz__9_14_inner_macOut_2 = (($signed(_zz__9_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_14_inner_activation;
    end else begin
      io_macOut = _9_14_inner_macOut;
    end
  end

  assign _zz__9_14_inner_macOut = ($signed(_zz__zz__9_14_inner_macOut) + $signed(_zz__zz__9_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_14_inner_activation <= 8'h00;
      _9_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_14_inner_activation <= io_addInput;
      end else begin
        _9_14_inner_macOut <= _zz__9_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_301 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_13_inner_macOut;
  wire       [15:0]   _zz__zz__9_13_inner_macOut_1;
  wire       [15:0]   _zz__9_13_inner_macOut_1;
  wire       [15:0]   _zz__9_13_inner_macOut_2;
  reg        [7:0]    _9_13_inner_activation;
  reg        [7:0]    _9_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_13_inner_macOut;

  assign _zz__zz__9_13_inner_macOut = ($signed(io_mulInput) * $signed(_9_13_inner_activation));
  assign _zz__zz__9_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_13_inner_macOut)) ? 16'h007f : _zz__9_13_inner_macOut_2);
  assign _zz__9_13_inner_macOut_2 = (($signed(_zz__9_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_13_inner_activation;
    end else begin
      io_macOut = _9_13_inner_macOut;
    end
  end

  assign _zz__9_13_inner_macOut = ($signed(_zz__zz__9_13_inner_macOut) + $signed(_zz__zz__9_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_13_inner_activation <= 8'h00;
      _9_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_13_inner_activation <= io_addInput;
      end else begin
        _9_13_inner_macOut <= _zz__9_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_300 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_12_inner_macOut;
  wire       [15:0]   _zz__zz__9_12_inner_macOut_1;
  wire       [15:0]   _zz__9_12_inner_macOut_1;
  wire       [15:0]   _zz__9_12_inner_macOut_2;
  reg        [7:0]    _9_12_inner_activation;
  reg        [7:0]    _9_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_12_inner_macOut;

  assign _zz__zz__9_12_inner_macOut = ($signed(io_mulInput) * $signed(_9_12_inner_activation));
  assign _zz__zz__9_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_12_inner_macOut)) ? 16'h007f : _zz__9_12_inner_macOut_2);
  assign _zz__9_12_inner_macOut_2 = (($signed(_zz__9_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_12_inner_activation;
    end else begin
      io_macOut = _9_12_inner_macOut;
    end
  end

  assign _zz__9_12_inner_macOut = ($signed(_zz__zz__9_12_inner_macOut) + $signed(_zz__zz__9_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_12_inner_activation <= 8'h00;
      _9_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_12_inner_activation <= io_addInput;
      end else begin
        _9_12_inner_macOut <= _zz__9_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_299 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_11_inner_macOut;
  wire       [15:0]   _zz__zz__9_11_inner_macOut_1;
  wire       [15:0]   _zz__9_11_inner_macOut_1;
  wire       [15:0]   _zz__9_11_inner_macOut_2;
  reg        [7:0]    _9_11_inner_activation;
  reg        [7:0]    _9_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_11_inner_macOut;

  assign _zz__zz__9_11_inner_macOut = ($signed(io_mulInput) * $signed(_9_11_inner_activation));
  assign _zz__zz__9_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_11_inner_macOut)) ? 16'h007f : _zz__9_11_inner_macOut_2);
  assign _zz__9_11_inner_macOut_2 = (($signed(_zz__9_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_11_inner_activation;
    end else begin
      io_macOut = _9_11_inner_macOut;
    end
  end

  assign _zz__9_11_inner_macOut = ($signed(_zz__zz__9_11_inner_macOut) + $signed(_zz__zz__9_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_11_inner_activation <= 8'h00;
      _9_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_11_inner_activation <= io_addInput;
      end else begin
        _9_11_inner_macOut <= _zz__9_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_298 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_10_inner_macOut;
  wire       [15:0]   _zz__zz__9_10_inner_macOut_1;
  wire       [15:0]   _zz__9_10_inner_macOut_1;
  wire       [15:0]   _zz__9_10_inner_macOut_2;
  reg        [7:0]    _9_10_inner_activation;
  reg        [7:0]    _9_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_10_inner_macOut;

  assign _zz__zz__9_10_inner_macOut = ($signed(io_mulInput) * $signed(_9_10_inner_activation));
  assign _zz__zz__9_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_10_inner_macOut)) ? 16'h007f : _zz__9_10_inner_macOut_2);
  assign _zz__9_10_inner_macOut_2 = (($signed(_zz__9_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_10_inner_activation;
    end else begin
      io_macOut = _9_10_inner_macOut;
    end
  end

  assign _zz__9_10_inner_macOut = ($signed(_zz__zz__9_10_inner_macOut) + $signed(_zz__zz__9_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_10_inner_activation <= 8'h00;
      _9_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_10_inner_activation <= io_addInput;
      end else begin
        _9_10_inner_macOut <= _zz__9_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_297 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_9_inner_macOut;
  wire       [15:0]   _zz__zz__9_9_inner_macOut_1;
  wire       [15:0]   _zz__9_9_inner_macOut_1;
  wire       [15:0]   _zz__9_9_inner_macOut_2;
  reg        [7:0]    _9_9_inner_activation;
  reg        [7:0]    _9_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_9_inner_macOut;

  assign _zz__zz__9_9_inner_macOut = ($signed(io_mulInput) * $signed(_9_9_inner_activation));
  assign _zz__zz__9_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_9_inner_macOut)) ? 16'h007f : _zz__9_9_inner_macOut_2);
  assign _zz__9_9_inner_macOut_2 = (($signed(_zz__9_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_9_inner_activation;
    end else begin
      io_macOut = _9_9_inner_macOut;
    end
  end

  assign _zz__9_9_inner_macOut = ($signed(_zz__zz__9_9_inner_macOut) + $signed(_zz__zz__9_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_9_inner_activation <= 8'h00;
      _9_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_9_inner_activation <= io_addInput;
      end else begin
        _9_9_inner_macOut <= _zz__9_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_296 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_8_inner_macOut;
  wire       [15:0]   _zz__zz__9_8_inner_macOut_1;
  wire       [15:0]   _zz__9_8_inner_macOut_1;
  wire       [15:0]   _zz__9_8_inner_macOut_2;
  reg        [7:0]    _9_8_inner_activation;
  reg        [7:0]    _9_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_8_inner_macOut;

  assign _zz__zz__9_8_inner_macOut = ($signed(io_mulInput) * $signed(_9_8_inner_activation));
  assign _zz__zz__9_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_8_inner_macOut)) ? 16'h007f : _zz__9_8_inner_macOut_2);
  assign _zz__9_8_inner_macOut_2 = (($signed(_zz__9_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_8_inner_activation;
    end else begin
      io_macOut = _9_8_inner_macOut;
    end
  end

  assign _zz__9_8_inner_macOut = ($signed(_zz__zz__9_8_inner_macOut) + $signed(_zz__zz__9_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_8_inner_activation <= 8'h00;
      _9_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_8_inner_activation <= io_addInput;
      end else begin
        _9_8_inner_macOut <= _zz__9_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_295 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_7_inner_macOut;
  wire       [15:0]   _zz__zz__9_7_inner_macOut_1;
  wire       [15:0]   _zz__9_7_inner_macOut_1;
  wire       [15:0]   _zz__9_7_inner_macOut_2;
  reg        [7:0]    _9_7_inner_activation;
  reg        [7:0]    _9_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_7_inner_macOut;

  assign _zz__zz__9_7_inner_macOut = ($signed(io_mulInput) * $signed(_9_7_inner_activation));
  assign _zz__zz__9_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_7_inner_macOut)) ? 16'h007f : _zz__9_7_inner_macOut_2);
  assign _zz__9_7_inner_macOut_2 = (($signed(_zz__9_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_7_inner_activation;
    end else begin
      io_macOut = _9_7_inner_macOut;
    end
  end

  assign _zz__9_7_inner_macOut = ($signed(_zz__zz__9_7_inner_macOut) + $signed(_zz__zz__9_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_7_inner_activation <= 8'h00;
      _9_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_7_inner_activation <= io_addInput;
      end else begin
        _9_7_inner_macOut <= _zz__9_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_294 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_6_inner_macOut;
  wire       [15:0]   _zz__zz__9_6_inner_macOut_1;
  wire       [15:0]   _zz__9_6_inner_macOut_1;
  wire       [15:0]   _zz__9_6_inner_macOut_2;
  reg        [7:0]    _9_6_inner_activation;
  reg        [7:0]    _9_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_6_inner_macOut;

  assign _zz__zz__9_6_inner_macOut = ($signed(io_mulInput) * $signed(_9_6_inner_activation));
  assign _zz__zz__9_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_6_inner_macOut)) ? 16'h007f : _zz__9_6_inner_macOut_2);
  assign _zz__9_6_inner_macOut_2 = (($signed(_zz__9_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_6_inner_activation;
    end else begin
      io_macOut = _9_6_inner_macOut;
    end
  end

  assign _zz__9_6_inner_macOut = ($signed(_zz__zz__9_6_inner_macOut) + $signed(_zz__zz__9_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_6_inner_activation <= 8'h00;
      _9_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_6_inner_activation <= io_addInput;
      end else begin
        _9_6_inner_macOut <= _zz__9_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_293 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_5_inner_macOut;
  wire       [15:0]   _zz__zz__9_5_inner_macOut_1;
  wire       [15:0]   _zz__9_5_inner_macOut_1;
  wire       [15:0]   _zz__9_5_inner_macOut_2;
  reg        [7:0]    _9_5_inner_activation;
  reg        [7:0]    _9_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_5_inner_macOut;

  assign _zz__zz__9_5_inner_macOut = ($signed(io_mulInput) * $signed(_9_5_inner_activation));
  assign _zz__zz__9_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_5_inner_macOut)) ? 16'h007f : _zz__9_5_inner_macOut_2);
  assign _zz__9_5_inner_macOut_2 = (($signed(_zz__9_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_5_inner_activation;
    end else begin
      io_macOut = _9_5_inner_macOut;
    end
  end

  assign _zz__9_5_inner_macOut = ($signed(_zz__zz__9_5_inner_macOut) + $signed(_zz__zz__9_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_5_inner_activation <= 8'h00;
      _9_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_5_inner_activation <= io_addInput;
      end else begin
        _9_5_inner_macOut <= _zz__9_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_292 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_4_inner_macOut;
  wire       [15:0]   _zz__zz__9_4_inner_macOut_1;
  wire       [15:0]   _zz__9_4_inner_macOut_1;
  wire       [15:0]   _zz__9_4_inner_macOut_2;
  reg        [7:0]    _9_4_inner_activation;
  reg        [7:0]    _9_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_4_inner_macOut;

  assign _zz__zz__9_4_inner_macOut = ($signed(io_mulInput) * $signed(_9_4_inner_activation));
  assign _zz__zz__9_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_4_inner_macOut)) ? 16'h007f : _zz__9_4_inner_macOut_2);
  assign _zz__9_4_inner_macOut_2 = (($signed(_zz__9_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_4_inner_activation;
    end else begin
      io_macOut = _9_4_inner_macOut;
    end
  end

  assign _zz__9_4_inner_macOut = ($signed(_zz__zz__9_4_inner_macOut) + $signed(_zz__zz__9_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_4_inner_activation <= 8'h00;
      _9_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_4_inner_activation <= io_addInput;
      end else begin
        _9_4_inner_macOut <= _zz__9_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_291 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_3_inner_macOut;
  wire       [15:0]   _zz__zz__9_3_inner_macOut_1;
  wire       [15:0]   _zz__9_3_inner_macOut_1;
  wire       [15:0]   _zz__9_3_inner_macOut_2;
  reg        [7:0]    _9_3_inner_activation;
  reg        [7:0]    _9_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_3_inner_macOut;

  assign _zz__zz__9_3_inner_macOut = ($signed(io_mulInput) * $signed(_9_3_inner_activation));
  assign _zz__zz__9_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_3_inner_macOut)) ? 16'h007f : _zz__9_3_inner_macOut_2);
  assign _zz__9_3_inner_macOut_2 = (($signed(_zz__9_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_3_inner_activation;
    end else begin
      io_macOut = _9_3_inner_macOut;
    end
  end

  assign _zz__9_3_inner_macOut = ($signed(_zz__zz__9_3_inner_macOut) + $signed(_zz__zz__9_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_3_inner_activation <= 8'h00;
      _9_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_3_inner_activation <= io_addInput;
      end else begin
        _9_3_inner_macOut <= _zz__9_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_290 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_2_inner_macOut;
  wire       [15:0]   _zz__zz__9_2_inner_macOut_1;
  wire       [15:0]   _zz__9_2_inner_macOut_1;
  wire       [15:0]   _zz__9_2_inner_macOut_2;
  reg        [7:0]    _9_2_inner_activation;
  reg        [7:0]    _9_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_2_inner_macOut;

  assign _zz__zz__9_2_inner_macOut = ($signed(io_mulInput) * $signed(_9_2_inner_activation));
  assign _zz__zz__9_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_2_inner_macOut)) ? 16'h007f : _zz__9_2_inner_macOut_2);
  assign _zz__9_2_inner_macOut_2 = (($signed(_zz__9_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_2_inner_activation;
    end else begin
      io_macOut = _9_2_inner_macOut;
    end
  end

  assign _zz__9_2_inner_macOut = ($signed(_zz__zz__9_2_inner_macOut) + $signed(_zz__zz__9_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_2_inner_activation <= 8'h00;
      _9_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_2_inner_activation <= io_addInput;
      end else begin
        _9_2_inner_macOut <= _zz__9_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_289 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_1_inner_macOut;
  wire       [15:0]   _zz__zz__9_1_inner_macOut_1;
  wire       [15:0]   _zz__9_1_inner_macOut_1;
  wire       [15:0]   _zz__9_1_inner_macOut_2;
  reg        [7:0]    _9_1_inner_activation;
  reg        [7:0]    _9_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_1_inner_macOut;

  assign _zz__zz__9_1_inner_macOut = ($signed(io_mulInput) * $signed(_9_1_inner_activation));
  assign _zz__zz__9_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_1_inner_macOut)) ? 16'h007f : _zz__9_1_inner_macOut_2);
  assign _zz__9_1_inner_macOut_2 = (($signed(_zz__9_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_1_inner_activation;
    end else begin
      io_macOut = _9_1_inner_macOut;
    end
  end

  assign _zz__9_1_inner_macOut = ($signed(_zz__zz__9_1_inner_macOut) + $signed(_zz__zz__9_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_1_inner_activation <= 8'h00;
      _9_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_1_inner_activation <= io_addInput;
      end else begin
        _9_1_inner_macOut <= _zz__9_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_288 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__9_0_inner_macOut;
  wire       [15:0]   _zz__zz__9_0_inner_macOut_1;
  wire       [15:0]   _zz__9_0_inner_macOut_1;
  wire       [15:0]   _zz__9_0_inner_macOut_2;
  reg        [7:0]    _9_0_inner_activation;
  reg        [7:0]    _9_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__9_0_inner_macOut;

  assign _zz__zz__9_0_inner_macOut = ($signed(io_mulInput) * $signed(_9_0_inner_activation));
  assign _zz__zz__9_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__9_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__9_0_inner_macOut)) ? 16'h007f : _zz__9_0_inner_macOut_2);
  assign _zz__9_0_inner_macOut_2 = (($signed(_zz__9_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__9_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _9_0_inner_activation;
    end else begin
      io_macOut = _9_0_inner_macOut;
    end
  end

  assign _zz__9_0_inner_macOut = ($signed(_zz__zz__9_0_inner_macOut) + $signed(_zz__zz__9_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _9_0_inner_activation <= 8'h00;
      _9_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _9_0_inner_activation <= io_addInput;
      end else begin
        _9_0_inner_macOut <= _zz__9_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_287 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_31_inner_macOut;
  wire       [15:0]   _zz__zz__8_31_inner_macOut_1;
  wire       [15:0]   _zz__8_31_inner_macOut_1;
  wire       [15:0]   _zz__8_31_inner_macOut_2;
  reg        [7:0]    _8_31_inner_activation;
  reg        [7:0]    _8_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_31_inner_macOut;

  assign _zz__zz__8_31_inner_macOut = ($signed(io_mulInput) * $signed(_8_31_inner_activation));
  assign _zz__zz__8_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_31_inner_macOut)) ? 16'h007f : _zz__8_31_inner_macOut_2);
  assign _zz__8_31_inner_macOut_2 = (($signed(_zz__8_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_31_inner_activation;
    end else begin
      io_macOut = _8_31_inner_macOut;
    end
  end

  assign _zz__8_31_inner_macOut = ($signed(_zz__zz__8_31_inner_macOut) + $signed(_zz__zz__8_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_31_inner_activation <= 8'h00;
      _8_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_31_inner_activation <= io_addInput;
      end else begin
        _8_31_inner_macOut <= _zz__8_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_286 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_30_inner_macOut;
  wire       [15:0]   _zz__zz__8_30_inner_macOut_1;
  wire       [15:0]   _zz__8_30_inner_macOut_1;
  wire       [15:0]   _zz__8_30_inner_macOut_2;
  reg        [7:0]    _8_30_inner_activation;
  reg        [7:0]    _8_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_30_inner_macOut;

  assign _zz__zz__8_30_inner_macOut = ($signed(io_mulInput) * $signed(_8_30_inner_activation));
  assign _zz__zz__8_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_30_inner_macOut)) ? 16'h007f : _zz__8_30_inner_macOut_2);
  assign _zz__8_30_inner_macOut_2 = (($signed(_zz__8_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_30_inner_activation;
    end else begin
      io_macOut = _8_30_inner_macOut;
    end
  end

  assign _zz__8_30_inner_macOut = ($signed(_zz__zz__8_30_inner_macOut) + $signed(_zz__zz__8_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_30_inner_activation <= 8'h00;
      _8_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_30_inner_activation <= io_addInput;
      end else begin
        _8_30_inner_macOut <= _zz__8_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_285 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_29_inner_macOut;
  wire       [15:0]   _zz__zz__8_29_inner_macOut_1;
  wire       [15:0]   _zz__8_29_inner_macOut_1;
  wire       [15:0]   _zz__8_29_inner_macOut_2;
  reg        [7:0]    _8_29_inner_activation;
  reg        [7:0]    _8_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_29_inner_macOut;

  assign _zz__zz__8_29_inner_macOut = ($signed(io_mulInput) * $signed(_8_29_inner_activation));
  assign _zz__zz__8_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_29_inner_macOut)) ? 16'h007f : _zz__8_29_inner_macOut_2);
  assign _zz__8_29_inner_macOut_2 = (($signed(_zz__8_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_29_inner_activation;
    end else begin
      io_macOut = _8_29_inner_macOut;
    end
  end

  assign _zz__8_29_inner_macOut = ($signed(_zz__zz__8_29_inner_macOut) + $signed(_zz__zz__8_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_29_inner_activation <= 8'h00;
      _8_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_29_inner_activation <= io_addInput;
      end else begin
        _8_29_inner_macOut <= _zz__8_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_284 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_28_inner_macOut;
  wire       [15:0]   _zz__zz__8_28_inner_macOut_1;
  wire       [15:0]   _zz__8_28_inner_macOut_1;
  wire       [15:0]   _zz__8_28_inner_macOut_2;
  reg        [7:0]    _8_28_inner_activation;
  reg        [7:0]    _8_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_28_inner_macOut;

  assign _zz__zz__8_28_inner_macOut = ($signed(io_mulInput) * $signed(_8_28_inner_activation));
  assign _zz__zz__8_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_28_inner_macOut)) ? 16'h007f : _zz__8_28_inner_macOut_2);
  assign _zz__8_28_inner_macOut_2 = (($signed(_zz__8_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_28_inner_activation;
    end else begin
      io_macOut = _8_28_inner_macOut;
    end
  end

  assign _zz__8_28_inner_macOut = ($signed(_zz__zz__8_28_inner_macOut) + $signed(_zz__zz__8_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_28_inner_activation <= 8'h00;
      _8_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_28_inner_activation <= io_addInput;
      end else begin
        _8_28_inner_macOut <= _zz__8_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_283 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_27_inner_macOut;
  wire       [15:0]   _zz__zz__8_27_inner_macOut_1;
  wire       [15:0]   _zz__8_27_inner_macOut_1;
  wire       [15:0]   _zz__8_27_inner_macOut_2;
  reg        [7:0]    _8_27_inner_activation;
  reg        [7:0]    _8_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_27_inner_macOut;

  assign _zz__zz__8_27_inner_macOut = ($signed(io_mulInput) * $signed(_8_27_inner_activation));
  assign _zz__zz__8_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_27_inner_macOut)) ? 16'h007f : _zz__8_27_inner_macOut_2);
  assign _zz__8_27_inner_macOut_2 = (($signed(_zz__8_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_27_inner_activation;
    end else begin
      io_macOut = _8_27_inner_macOut;
    end
  end

  assign _zz__8_27_inner_macOut = ($signed(_zz__zz__8_27_inner_macOut) + $signed(_zz__zz__8_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_27_inner_activation <= 8'h00;
      _8_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_27_inner_activation <= io_addInput;
      end else begin
        _8_27_inner_macOut <= _zz__8_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_282 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_26_inner_macOut;
  wire       [15:0]   _zz__zz__8_26_inner_macOut_1;
  wire       [15:0]   _zz__8_26_inner_macOut_1;
  wire       [15:0]   _zz__8_26_inner_macOut_2;
  reg        [7:0]    _8_26_inner_activation;
  reg        [7:0]    _8_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_26_inner_macOut;

  assign _zz__zz__8_26_inner_macOut = ($signed(io_mulInput) * $signed(_8_26_inner_activation));
  assign _zz__zz__8_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_26_inner_macOut)) ? 16'h007f : _zz__8_26_inner_macOut_2);
  assign _zz__8_26_inner_macOut_2 = (($signed(_zz__8_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_26_inner_activation;
    end else begin
      io_macOut = _8_26_inner_macOut;
    end
  end

  assign _zz__8_26_inner_macOut = ($signed(_zz__zz__8_26_inner_macOut) + $signed(_zz__zz__8_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_26_inner_activation <= 8'h00;
      _8_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_26_inner_activation <= io_addInput;
      end else begin
        _8_26_inner_macOut <= _zz__8_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_281 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_25_inner_macOut;
  wire       [15:0]   _zz__zz__8_25_inner_macOut_1;
  wire       [15:0]   _zz__8_25_inner_macOut_1;
  wire       [15:0]   _zz__8_25_inner_macOut_2;
  reg        [7:0]    _8_25_inner_activation;
  reg        [7:0]    _8_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_25_inner_macOut;

  assign _zz__zz__8_25_inner_macOut = ($signed(io_mulInput) * $signed(_8_25_inner_activation));
  assign _zz__zz__8_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_25_inner_macOut)) ? 16'h007f : _zz__8_25_inner_macOut_2);
  assign _zz__8_25_inner_macOut_2 = (($signed(_zz__8_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_25_inner_activation;
    end else begin
      io_macOut = _8_25_inner_macOut;
    end
  end

  assign _zz__8_25_inner_macOut = ($signed(_zz__zz__8_25_inner_macOut) + $signed(_zz__zz__8_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_25_inner_activation <= 8'h00;
      _8_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_25_inner_activation <= io_addInput;
      end else begin
        _8_25_inner_macOut <= _zz__8_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_280 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_24_inner_macOut;
  wire       [15:0]   _zz__zz__8_24_inner_macOut_1;
  wire       [15:0]   _zz__8_24_inner_macOut_1;
  wire       [15:0]   _zz__8_24_inner_macOut_2;
  reg        [7:0]    _8_24_inner_activation;
  reg        [7:0]    _8_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_24_inner_macOut;

  assign _zz__zz__8_24_inner_macOut = ($signed(io_mulInput) * $signed(_8_24_inner_activation));
  assign _zz__zz__8_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_24_inner_macOut)) ? 16'h007f : _zz__8_24_inner_macOut_2);
  assign _zz__8_24_inner_macOut_2 = (($signed(_zz__8_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_24_inner_activation;
    end else begin
      io_macOut = _8_24_inner_macOut;
    end
  end

  assign _zz__8_24_inner_macOut = ($signed(_zz__zz__8_24_inner_macOut) + $signed(_zz__zz__8_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_24_inner_activation <= 8'h00;
      _8_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_24_inner_activation <= io_addInput;
      end else begin
        _8_24_inner_macOut <= _zz__8_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_279 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_23_inner_macOut;
  wire       [15:0]   _zz__zz__8_23_inner_macOut_1;
  wire       [15:0]   _zz__8_23_inner_macOut_1;
  wire       [15:0]   _zz__8_23_inner_macOut_2;
  reg        [7:0]    _8_23_inner_activation;
  reg        [7:0]    _8_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_23_inner_macOut;

  assign _zz__zz__8_23_inner_macOut = ($signed(io_mulInput) * $signed(_8_23_inner_activation));
  assign _zz__zz__8_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_23_inner_macOut)) ? 16'h007f : _zz__8_23_inner_macOut_2);
  assign _zz__8_23_inner_macOut_2 = (($signed(_zz__8_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_23_inner_activation;
    end else begin
      io_macOut = _8_23_inner_macOut;
    end
  end

  assign _zz__8_23_inner_macOut = ($signed(_zz__zz__8_23_inner_macOut) + $signed(_zz__zz__8_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_23_inner_activation <= 8'h00;
      _8_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_23_inner_activation <= io_addInput;
      end else begin
        _8_23_inner_macOut <= _zz__8_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_278 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_22_inner_macOut;
  wire       [15:0]   _zz__zz__8_22_inner_macOut_1;
  wire       [15:0]   _zz__8_22_inner_macOut_1;
  wire       [15:0]   _zz__8_22_inner_macOut_2;
  reg        [7:0]    _8_22_inner_activation;
  reg        [7:0]    _8_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_22_inner_macOut;

  assign _zz__zz__8_22_inner_macOut = ($signed(io_mulInput) * $signed(_8_22_inner_activation));
  assign _zz__zz__8_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_22_inner_macOut)) ? 16'h007f : _zz__8_22_inner_macOut_2);
  assign _zz__8_22_inner_macOut_2 = (($signed(_zz__8_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_22_inner_activation;
    end else begin
      io_macOut = _8_22_inner_macOut;
    end
  end

  assign _zz__8_22_inner_macOut = ($signed(_zz__zz__8_22_inner_macOut) + $signed(_zz__zz__8_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_22_inner_activation <= 8'h00;
      _8_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_22_inner_activation <= io_addInput;
      end else begin
        _8_22_inner_macOut <= _zz__8_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_277 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_21_inner_macOut;
  wire       [15:0]   _zz__zz__8_21_inner_macOut_1;
  wire       [15:0]   _zz__8_21_inner_macOut_1;
  wire       [15:0]   _zz__8_21_inner_macOut_2;
  reg        [7:0]    _8_21_inner_activation;
  reg        [7:0]    _8_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_21_inner_macOut;

  assign _zz__zz__8_21_inner_macOut = ($signed(io_mulInput) * $signed(_8_21_inner_activation));
  assign _zz__zz__8_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_21_inner_macOut)) ? 16'h007f : _zz__8_21_inner_macOut_2);
  assign _zz__8_21_inner_macOut_2 = (($signed(_zz__8_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_21_inner_activation;
    end else begin
      io_macOut = _8_21_inner_macOut;
    end
  end

  assign _zz__8_21_inner_macOut = ($signed(_zz__zz__8_21_inner_macOut) + $signed(_zz__zz__8_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_21_inner_activation <= 8'h00;
      _8_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_21_inner_activation <= io_addInput;
      end else begin
        _8_21_inner_macOut <= _zz__8_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_276 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_20_inner_macOut;
  wire       [15:0]   _zz__zz__8_20_inner_macOut_1;
  wire       [15:0]   _zz__8_20_inner_macOut_1;
  wire       [15:0]   _zz__8_20_inner_macOut_2;
  reg        [7:0]    _8_20_inner_activation;
  reg        [7:0]    _8_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_20_inner_macOut;

  assign _zz__zz__8_20_inner_macOut = ($signed(io_mulInput) * $signed(_8_20_inner_activation));
  assign _zz__zz__8_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_20_inner_macOut)) ? 16'h007f : _zz__8_20_inner_macOut_2);
  assign _zz__8_20_inner_macOut_2 = (($signed(_zz__8_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_20_inner_activation;
    end else begin
      io_macOut = _8_20_inner_macOut;
    end
  end

  assign _zz__8_20_inner_macOut = ($signed(_zz__zz__8_20_inner_macOut) + $signed(_zz__zz__8_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_20_inner_activation <= 8'h00;
      _8_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_20_inner_activation <= io_addInput;
      end else begin
        _8_20_inner_macOut <= _zz__8_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_275 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_19_inner_macOut;
  wire       [15:0]   _zz__zz__8_19_inner_macOut_1;
  wire       [15:0]   _zz__8_19_inner_macOut_1;
  wire       [15:0]   _zz__8_19_inner_macOut_2;
  reg        [7:0]    _8_19_inner_activation;
  reg        [7:0]    _8_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_19_inner_macOut;

  assign _zz__zz__8_19_inner_macOut = ($signed(io_mulInput) * $signed(_8_19_inner_activation));
  assign _zz__zz__8_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_19_inner_macOut)) ? 16'h007f : _zz__8_19_inner_macOut_2);
  assign _zz__8_19_inner_macOut_2 = (($signed(_zz__8_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_19_inner_activation;
    end else begin
      io_macOut = _8_19_inner_macOut;
    end
  end

  assign _zz__8_19_inner_macOut = ($signed(_zz__zz__8_19_inner_macOut) + $signed(_zz__zz__8_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_19_inner_activation <= 8'h00;
      _8_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_19_inner_activation <= io_addInput;
      end else begin
        _8_19_inner_macOut <= _zz__8_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_274 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_18_inner_macOut;
  wire       [15:0]   _zz__zz__8_18_inner_macOut_1;
  wire       [15:0]   _zz__8_18_inner_macOut_1;
  wire       [15:0]   _zz__8_18_inner_macOut_2;
  reg        [7:0]    _8_18_inner_activation;
  reg        [7:0]    _8_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_18_inner_macOut;

  assign _zz__zz__8_18_inner_macOut = ($signed(io_mulInput) * $signed(_8_18_inner_activation));
  assign _zz__zz__8_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_18_inner_macOut)) ? 16'h007f : _zz__8_18_inner_macOut_2);
  assign _zz__8_18_inner_macOut_2 = (($signed(_zz__8_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_18_inner_activation;
    end else begin
      io_macOut = _8_18_inner_macOut;
    end
  end

  assign _zz__8_18_inner_macOut = ($signed(_zz__zz__8_18_inner_macOut) + $signed(_zz__zz__8_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_18_inner_activation <= 8'h00;
      _8_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_18_inner_activation <= io_addInput;
      end else begin
        _8_18_inner_macOut <= _zz__8_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_273 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_17_inner_macOut;
  wire       [15:0]   _zz__zz__8_17_inner_macOut_1;
  wire       [15:0]   _zz__8_17_inner_macOut_1;
  wire       [15:0]   _zz__8_17_inner_macOut_2;
  reg        [7:0]    _8_17_inner_activation;
  reg        [7:0]    _8_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_17_inner_macOut;

  assign _zz__zz__8_17_inner_macOut = ($signed(io_mulInput) * $signed(_8_17_inner_activation));
  assign _zz__zz__8_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_17_inner_macOut)) ? 16'h007f : _zz__8_17_inner_macOut_2);
  assign _zz__8_17_inner_macOut_2 = (($signed(_zz__8_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_17_inner_activation;
    end else begin
      io_macOut = _8_17_inner_macOut;
    end
  end

  assign _zz__8_17_inner_macOut = ($signed(_zz__zz__8_17_inner_macOut) + $signed(_zz__zz__8_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_17_inner_activation <= 8'h00;
      _8_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_17_inner_activation <= io_addInput;
      end else begin
        _8_17_inner_macOut <= _zz__8_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_272 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_16_inner_macOut;
  wire       [15:0]   _zz__zz__8_16_inner_macOut_1;
  wire       [15:0]   _zz__8_16_inner_macOut_1;
  wire       [15:0]   _zz__8_16_inner_macOut_2;
  reg        [7:0]    _8_16_inner_activation;
  reg        [7:0]    _8_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_16_inner_macOut;

  assign _zz__zz__8_16_inner_macOut = ($signed(io_mulInput) * $signed(_8_16_inner_activation));
  assign _zz__zz__8_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_16_inner_macOut)) ? 16'h007f : _zz__8_16_inner_macOut_2);
  assign _zz__8_16_inner_macOut_2 = (($signed(_zz__8_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_16_inner_activation;
    end else begin
      io_macOut = _8_16_inner_macOut;
    end
  end

  assign _zz__8_16_inner_macOut = ($signed(_zz__zz__8_16_inner_macOut) + $signed(_zz__zz__8_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_16_inner_activation <= 8'h00;
      _8_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_16_inner_activation <= io_addInput;
      end else begin
        _8_16_inner_macOut <= _zz__8_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_271 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_15_inner_macOut;
  wire       [15:0]   _zz__zz__8_15_inner_macOut_1;
  wire       [15:0]   _zz__8_15_inner_macOut_1;
  wire       [15:0]   _zz__8_15_inner_macOut_2;
  reg        [7:0]    _8_15_inner_activation;
  reg        [7:0]    _8_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_15_inner_macOut;

  assign _zz__zz__8_15_inner_macOut = ($signed(io_mulInput) * $signed(_8_15_inner_activation));
  assign _zz__zz__8_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_15_inner_macOut)) ? 16'h007f : _zz__8_15_inner_macOut_2);
  assign _zz__8_15_inner_macOut_2 = (($signed(_zz__8_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_15_inner_activation;
    end else begin
      io_macOut = _8_15_inner_macOut;
    end
  end

  assign _zz__8_15_inner_macOut = ($signed(_zz__zz__8_15_inner_macOut) + $signed(_zz__zz__8_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_15_inner_activation <= 8'h00;
      _8_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_15_inner_activation <= io_addInput;
      end else begin
        _8_15_inner_macOut <= _zz__8_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_270 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_14_inner_macOut;
  wire       [15:0]   _zz__zz__8_14_inner_macOut_1;
  wire       [15:0]   _zz__8_14_inner_macOut_1;
  wire       [15:0]   _zz__8_14_inner_macOut_2;
  reg        [7:0]    _8_14_inner_activation;
  reg        [7:0]    _8_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_14_inner_macOut;

  assign _zz__zz__8_14_inner_macOut = ($signed(io_mulInput) * $signed(_8_14_inner_activation));
  assign _zz__zz__8_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_14_inner_macOut)) ? 16'h007f : _zz__8_14_inner_macOut_2);
  assign _zz__8_14_inner_macOut_2 = (($signed(_zz__8_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_14_inner_activation;
    end else begin
      io_macOut = _8_14_inner_macOut;
    end
  end

  assign _zz__8_14_inner_macOut = ($signed(_zz__zz__8_14_inner_macOut) + $signed(_zz__zz__8_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_14_inner_activation <= 8'h00;
      _8_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_14_inner_activation <= io_addInput;
      end else begin
        _8_14_inner_macOut <= _zz__8_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_269 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_13_inner_macOut;
  wire       [15:0]   _zz__zz__8_13_inner_macOut_1;
  wire       [15:0]   _zz__8_13_inner_macOut_1;
  wire       [15:0]   _zz__8_13_inner_macOut_2;
  reg        [7:0]    _8_13_inner_activation;
  reg        [7:0]    _8_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_13_inner_macOut;

  assign _zz__zz__8_13_inner_macOut = ($signed(io_mulInput) * $signed(_8_13_inner_activation));
  assign _zz__zz__8_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_13_inner_macOut)) ? 16'h007f : _zz__8_13_inner_macOut_2);
  assign _zz__8_13_inner_macOut_2 = (($signed(_zz__8_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_13_inner_activation;
    end else begin
      io_macOut = _8_13_inner_macOut;
    end
  end

  assign _zz__8_13_inner_macOut = ($signed(_zz__zz__8_13_inner_macOut) + $signed(_zz__zz__8_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_13_inner_activation <= 8'h00;
      _8_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_13_inner_activation <= io_addInput;
      end else begin
        _8_13_inner_macOut <= _zz__8_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_268 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_12_inner_macOut;
  wire       [15:0]   _zz__zz__8_12_inner_macOut_1;
  wire       [15:0]   _zz__8_12_inner_macOut_1;
  wire       [15:0]   _zz__8_12_inner_macOut_2;
  reg        [7:0]    _8_12_inner_activation;
  reg        [7:0]    _8_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_12_inner_macOut;

  assign _zz__zz__8_12_inner_macOut = ($signed(io_mulInput) * $signed(_8_12_inner_activation));
  assign _zz__zz__8_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_12_inner_macOut)) ? 16'h007f : _zz__8_12_inner_macOut_2);
  assign _zz__8_12_inner_macOut_2 = (($signed(_zz__8_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_12_inner_activation;
    end else begin
      io_macOut = _8_12_inner_macOut;
    end
  end

  assign _zz__8_12_inner_macOut = ($signed(_zz__zz__8_12_inner_macOut) + $signed(_zz__zz__8_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_12_inner_activation <= 8'h00;
      _8_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_12_inner_activation <= io_addInput;
      end else begin
        _8_12_inner_macOut <= _zz__8_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_267 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_11_inner_macOut;
  wire       [15:0]   _zz__zz__8_11_inner_macOut_1;
  wire       [15:0]   _zz__8_11_inner_macOut_1;
  wire       [15:0]   _zz__8_11_inner_macOut_2;
  reg        [7:0]    _8_11_inner_activation;
  reg        [7:0]    _8_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_11_inner_macOut;

  assign _zz__zz__8_11_inner_macOut = ($signed(io_mulInput) * $signed(_8_11_inner_activation));
  assign _zz__zz__8_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_11_inner_macOut)) ? 16'h007f : _zz__8_11_inner_macOut_2);
  assign _zz__8_11_inner_macOut_2 = (($signed(_zz__8_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_11_inner_activation;
    end else begin
      io_macOut = _8_11_inner_macOut;
    end
  end

  assign _zz__8_11_inner_macOut = ($signed(_zz__zz__8_11_inner_macOut) + $signed(_zz__zz__8_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_11_inner_activation <= 8'h00;
      _8_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_11_inner_activation <= io_addInput;
      end else begin
        _8_11_inner_macOut <= _zz__8_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_266 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_10_inner_macOut;
  wire       [15:0]   _zz__zz__8_10_inner_macOut_1;
  wire       [15:0]   _zz__8_10_inner_macOut_1;
  wire       [15:0]   _zz__8_10_inner_macOut_2;
  reg        [7:0]    _8_10_inner_activation;
  reg        [7:0]    _8_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_10_inner_macOut;

  assign _zz__zz__8_10_inner_macOut = ($signed(io_mulInput) * $signed(_8_10_inner_activation));
  assign _zz__zz__8_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_10_inner_macOut)) ? 16'h007f : _zz__8_10_inner_macOut_2);
  assign _zz__8_10_inner_macOut_2 = (($signed(_zz__8_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_10_inner_activation;
    end else begin
      io_macOut = _8_10_inner_macOut;
    end
  end

  assign _zz__8_10_inner_macOut = ($signed(_zz__zz__8_10_inner_macOut) + $signed(_zz__zz__8_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_10_inner_activation <= 8'h00;
      _8_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_10_inner_activation <= io_addInput;
      end else begin
        _8_10_inner_macOut <= _zz__8_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_265 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_9_inner_macOut;
  wire       [15:0]   _zz__zz__8_9_inner_macOut_1;
  wire       [15:0]   _zz__8_9_inner_macOut_1;
  wire       [15:0]   _zz__8_9_inner_macOut_2;
  reg        [7:0]    _8_9_inner_activation;
  reg        [7:0]    _8_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_9_inner_macOut;

  assign _zz__zz__8_9_inner_macOut = ($signed(io_mulInput) * $signed(_8_9_inner_activation));
  assign _zz__zz__8_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_9_inner_macOut)) ? 16'h007f : _zz__8_9_inner_macOut_2);
  assign _zz__8_9_inner_macOut_2 = (($signed(_zz__8_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_9_inner_activation;
    end else begin
      io_macOut = _8_9_inner_macOut;
    end
  end

  assign _zz__8_9_inner_macOut = ($signed(_zz__zz__8_9_inner_macOut) + $signed(_zz__zz__8_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_9_inner_activation <= 8'h00;
      _8_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_9_inner_activation <= io_addInput;
      end else begin
        _8_9_inner_macOut <= _zz__8_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_264 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_8_inner_macOut;
  wire       [15:0]   _zz__zz__8_8_inner_macOut_1;
  wire       [15:0]   _zz__8_8_inner_macOut_1;
  wire       [15:0]   _zz__8_8_inner_macOut_2;
  reg        [7:0]    _8_8_inner_activation;
  reg        [7:0]    _8_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_8_inner_macOut;

  assign _zz__zz__8_8_inner_macOut = ($signed(io_mulInput) * $signed(_8_8_inner_activation));
  assign _zz__zz__8_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_8_inner_macOut)) ? 16'h007f : _zz__8_8_inner_macOut_2);
  assign _zz__8_8_inner_macOut_2 = (($signed(_zz__8_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_8_inner_activation;
    end else begin
      io_macOut = _8_8_inner_macOut;
    end
  end

  assign _zz__8_8_inner_macOut = ($signed(_zz__zz__8_8_inner_macOut) + $signed(_zz__zz__8_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_8_inner_activation <= 8'h00;
      _8_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_8_inner_activation <= io_addInput;
      end else begin
        _8_8_inner_macOut <= _zz__8_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_263 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_7_inner_macOut;
  wire       [15:0]   _zz__zz__8_7_inner_macOut_1;
  wire       [15:0]   _zz__8_7_inner_macOut_1;
  wire       [15:0]   _zz__8_7_inner_macOut_2;
  reg        [7:0]    _8_7_inner_activation;
  reg        [7:0]    _8_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_7_inner_macOut;

  assign _zz__zz__8_7_inner_macOut = ($signed(io_mulInput) * $signed(_8_7_inner_activation));
  assign _zz__zz__8_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_7_inner_macOut)) ? 16'h007f : _zz__8_7_inner_macOut_2);
  assign _zz__8_7_inner_macOut_2 = (($signed(_zz__8_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_7_inner_activation;
    end else begin
      io_macOut = _8_7_inner_macOut;
    end
  end

  assign _zz__8_7_inner_macOut = ($signed(_zz__zz__8_7_inner_macOut) + $signed(_zz__zz__8_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_7_inner_activation <= 8'h00;
      _8_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_7_inner_activation <= io_addInput;
      end else begin
        _8_7_inner_macOut <= _zz__8_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_262 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_6_inner_macOut;
  wire       [15:0]   _zz__zz__8_6_inner_macOut_1;
  wire       [15:0]   _zz__8_6_inner_macOut_1;
  wire       [15:0]   _zz__8_6_inner_macOut_2;
  reg        [7:0]    _8_6_inner_activation;
  reg        [7:0]    _8_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_6_inner_macOut;

  assign _zz__zz__8_6_inner_macOut = ($signed(io_mulInput) * $signed(_8_6_inner_activation));
  assign _zz__zz__8_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_6_inner_macOut)) ? 16'h007f : _zz__8_6_inner_macOut_2);
  assign _zz__8_6_inner_macOut_2 = (($signed(_zz__8_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_6_inner_activation;
    end else begin
      io_macOut = _8_6_inner_macOut;
    end
  end

  assign _zz__8_6_inner_macOut = ($signed(_zz__zz__8_6_inner_macOut) + $signed(_zz__zz__8_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_6_inner_activation <= 8'h00;
      _8_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_6_inner_activation <= io_addInput;
      end else begin
        _8_6_inner_macOut <= _zz__8_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_261 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_5_inner_macOut;
  wire       [15:0]   _zz__zz__8_5_inner_macOut_1;
  wire       [15:0]   _zz__8_5_inner_macOut_1;
  wire       [15:0]   _zz__8_5_inner_macOut_2;
  reg        [7:0]    _8_5_inner_activation;
  reg        [7:0]    _8_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_5_inner_macOut;

  assign _zz__zz__8_5_inner_macOut = ($signed(io_mulInput) * $signed(_8_5_inner_activation));
  assign _zz__zz__8_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_5_inner_macOut)) ? 16'h007f : _zz__8_5_inner_macOut_2);
  assign _zz__8_5_inner_macOut_2 = (($signed(_zz__8_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_5_inner_activation;
    end else begin
      io_macOut = _8_5_inner_macOut;
    end
  end

  assign _zz__8_5_inner_macOut = ($signed(_zz__zz__8_5_inner_macOut) + $signed(_zz__zz__8_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_5_inner_activation <= 8'h00;
      _8_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_5_inner_activation <= io_addInput;
      end else begin
        _8_5_inner_macOut <= _zz__8_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_260 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_4_inner_macOut;
  wire       [15:0]   _zz__zz__8_4_inner_macOut_1;
  wire       [15:0]   _zz__8_4_inner_macOut_1;
  wire       [15:0]   _zz__8_4_inner_macOut_2;
  reg        [7:0]    _8_4_inner_activation;
  reg        [7:0]    _8_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_4_inner_macOut;

  assign _zz__zz__8_4_inner_macOut = ($signed(io_mulInput) * $signed(_8_4_inner_activation));
  assign _zz__zz__8_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_4_inner_macOut)) ? 16'h007f : _zz__8_4_inner_macOut_2);
  assign _zz__8_4_inner_macOut_2 = (($signed(_zz__8_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_4_inner_activation;
    end else begin
      io_macOut = _8_4_inner_macOut;
    end
  end

  assign _zz__8_4_inner_macOut = ($signed(_zz__zz__8_4_inner_macOut) + $signed(_zz__zz__8_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_4_inner_activation <= 8'h00;
      _8_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_4_inner_activation <= io_addInput;
      end else begin
        _8_4_inner_macOut <= _zz__8_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_259 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_3_inner_macOut;
  wire       [15:0]   _zz__zz__8_3_inner_macOut_1;
  wire       [15:0]   _zz__8_3_inner_macOut_1;
  wire       [15:0]   _zz__8_3_inner_macOut_2;
  reg        [7:0]    _8_3_inner_activation;
  reg        [7:0]    _8_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_3_inner_macOut;

  assign _zz__zz__8_3_inner_macOut = ($signed(io_mulInput) * $signed(_8_3_inner_activation));
  assign _zz__zz__8_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_3_inner_macOut)) ? 16'h007f : _zz__8_3_inner_macOut_2);
  assign _zz__8_3_inner_macOut_2 = (($signed(_zz__8_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_3_inner_activation;
    end else begin
      io_macOut = _8_3_inner_macOut;
    end
  end

  assign _zz__8_3_inner_macOut = ($signed(_zz__zz__8_3_inner_macOut) + $signed(_zz__zz__8_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_3_inner_activation <= 8'h00;
      _8_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_3_inner_activation <= io_addInput;
      end else begin
        _8_3_inner_macOut <= _zz__8_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_258 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_2_inner_macOut;
  wire       [15:0]   _zz__zz__8_2_inner_macOut_1;
  wire       [15:0]   _zz__8_2_inner_macOut_1;
  wire       [15:0]   _zz__8_2_inner_macOut_2;
  reg        [7:0]    _8_2_inner_activation;
  reg        [7:0]    _8_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_2_inner_macOut;

  assign _zz__zz__8_2_inner_macOut = ($signed(io_mulInput) * $signed(_8_2_inner_activation));
  assign _zz__zz__8_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_2_inner_macOut)) ? 16'h007f : _zz__8_2_inner_macOut_2);
  assign _zz__8_2_inner_macOut_2 = (($signed(_zz__8_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_2_inner_activation;
    end else begin
      io_macOut = _8_2_inner_macOut;
    end
  end

  assign _zz__8_2_inner_macOut = ($signed(_zz__zz__8_2_inner_macOut) + $signed(_zz__zz__8_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_2_inner_activation <= 8'h00;
      _8_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_2_inner_activation <= io_addInput;
      end else begin
        _8_2_inner_macOut <= _zz__8_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_257 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_1_inner_macOut;
  wire       [15:0]   _zz__zz__8_1_inner_macOut_1;
  wire       [15:0]   _zz__8_1_inner_macOut_1;
  wire       [15:0]   _zz__8_1_inner_macOut_2;
  reg        [7:0]    _8_1_inner_activation;
  reg        [7:0]    _8_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_1_inner_macOut;

  assign _zz__zz__8_1_inner_macOut = ($signed(io_mulInput) * $signed(_8_1_inner_activation));
  assign _zz__zz__8_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_1_inner_macOut)) ? 16'h007f : _zz__8_1_inner_macOut_2);
  assign _zz__8_1_inner_macOut_2 = (($signed(_zz__8_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_1_inner_activation;
    end else begin
      io_macOut = _8_1_inner_macOut;
    end
  end

  assign _zz__8_1_inner_macOut = ($signed(_zz__zz__8_1_inner_macOut) + $signed(_zz__zz__8_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_1_inner_activation <= 8'h00;
      _8_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_1_inner_activation <= io_addInput;
      end else begin
        _8_1_inner_macOut <= _zz__8_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_256 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__8_0_inner_macOut;
  wire       [15:0]   _zz__zz__8_0_inner_macOut_1;
  wire       [15:0]   _zz__8_0_inner_macOut_1;
  wire       [15:0]   _zz__8_0_inner_macOut_2;
  reg        [7:0]    _8_0_inner_activation;
  reg        [7:0]    _8_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__8_0_inner_macOut;

  assign _zz__zz__8_0_inner_macOut = ($signed(io_mulInput) * $signed(_8_0_inner_activation));
  assign _zz__zz__8_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__8_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__8_0_inner_macOut)) ? 16'h007f : _zz__8_0_inner_macOut_2);
  assign _zz__8_0_inner_macOut_2 = (($signed(_zz__8_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__8_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _8_0_inner_activation;
    end else begin
      io_macOut = _8_0_inner_macOut;
    end
  end

  assign _zz__8_0_inner_macOut = ($signed(_zz__zz__8_0_inner_macOut) + $signed(_zz__zz__8_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _8_0_inner_activation <= 8'h00;
      _8_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _8_0_inner_activation <= io_addInput;
      end else begin
        _8_0_inner_macOut <= _zz__8_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_255 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_31_inner_macOut;
  wire       [15:0]   _zz__zz__7_31_inner_macOut_1;
  wire       [15:0]   _zz__7_31_inner_macOut_1;
  wire       [15:0]   _zz__7_31_inner_macOut_2;
  reg        [7:0]    _7_31_inner_activation;
  reg        [7:0]    _7_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_31_inner_macOut;

  assign _zz__zz__7_31_inner_macOut = ($signed(io_mulInput) * $signed(_7_31_inner_activation));
  assign _zz__zz__7_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_31_inner_macOut)) ? 16'h007f : _zz__7_31_inner_macOut_2);
  assign _zz__7_31_inner_macOut_2 = (($signed(_zz__7_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_31_inner_activation;
    end else begin
      io_macOut = _7_31_inner_macOut;
    end
  end

  assign _zz__7_31_inner_macOut = ($signed(_zz__zz__7_31_inner_macOut) + $signed(_zz__zz__7_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_31_inner_activation <= 8'h00;
      _7_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_31_inner_activation <= io_addInput;
      end else begin
        _7_31_inner_macOut <= _zz__7_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_254 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_30_inner_macOut;
  wire       [15:0]   _zz__zz__7_30_inner_macOut_1;
  wire       [15:0]   _zz__7_30_inner_macOut_1;
  wire       [15:0]   _zz__7_30_inner_macOut_2;
  reg        [7:0]    _7_30_inner_activation;
  reg        [7:0]    _7_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_30_inner_macOut;

  assign _zz__zz__7_30_inner_macOut = ($signed(io_mulInput) * $signed(_7_30_inner_activation));
  assign _zz__zz__7_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_30_inner_macOut)) ? 16'h007f : _zz__7_30_inner_macOut_2);
  assign _zz__7_30_inner_macOut_2 = (($signed(_zz__7_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_30_inner_activation;
    end else begin
      io_macOut = _7_30_inner_macOut;
    end
  end

  assign _zz__7_30_inner_macOut = ($signed(_zz__zz__7_30_inner_macOut) + $signed(_zz__zz__7_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_30_inner_activation <= 8'h00;
      _7_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_30_inner_activation <= io_addInput;
      end else begin
        _7_30_inner_macOut <= _zz__7_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_253 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_29_inner_macOut;
  wire       [15:0]   _zz__zz__7_29_inner_macOut_1;
  wire       [15:0]   _zz__7_29_inner_macOut_1;
  wire       [15:0]   _zz__7_29_inner_macOut_2;
  reg        [7:0]    _7_29_inner_activation;
  reg        [7:0]    _7_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_29_inner_macOut;

  assign _zz__zz__7_29_inner_macOut = ($signed(io_mulInput) * $signed(_7_29_inner_activation));
  assign _zz__zz__7_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_29_inner_macOut)) ? 16'h007f : _zz__7_29_inner_macOut_2);
  assign _zz__7_29_inner_macOut_2 = (($signed(_zz__7_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_29_inner_activation;
    end else begin
      io_macOut = _7_29_inner_macOut;
    end
  end

  assign _zz__7_29_inner_macOut = ($signed(_zz__zz__7_29_inner_macOut) + $signed(_zz__zz__7_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_29_inner_activation <= 8'h00;
      _7_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_29_inner_activation <= io_addInput;
      end else begin
        _7_29_inner_macOut <= _zz__7_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_252 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_28_inner_macOut;
  wire       [15:0]   _zz__zz__7_28_inner_macOut_1;
  wire       [15:0]   _zz__7_28_inner_macOut_1;
  wire       [15:0]   _zz__7_28_inner_macOut_2;
  reg        [7:0]    _7_28_inner_activation;
  reg        [7:0]    _7_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_28_inner_macOut;

  assign _zz__zz__7_28_inner_macOut = ($signed(io_mulInput) * $signed(_7_28_inner_activation));
  assign _zz__zz__7_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_28_inner_macOut)) ? 16'h007f : _zz__7_28_inner_macOut_2);
  assign _zz__7_28_inner_macOut_2 = (($signed(_zz__7_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_28_inner_activation;
    end else begin
      io_macOut = _7_28_inner_macOut;
    end
  end

  assign _zz__7_28_inner_macOut = ($signed(_zz__zz__7_28_inner_macOut) + $signed(_zz__zz__7_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_28_inner_activation <= 8'h00;
      _7_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_28_inner_activation <= io_addInput;
      end else begin
        _7_28_inner_macOut <= _zz__7_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_251 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_27_inner_macOut;
  wire       [15:0]   _zz__zz__7_27_inner_macOut_1;
  wire       [15:0]   _zz__7_27_inner_macOut_1;
  wire       [15:0]   _zz__7_27_inner_macOut_2;
  reg        [7:0]    _7_27_inner_activation;
  reg        [7:0]    _7_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_27_inner_macOut;

  assign _zz__zz__7_27_inner_macOut = ($signed(io_mulInput) * $signed(_7_27_inner_activation));
  assign _zz__zz__7_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_27_inner_macOut)) ? 16'h007f : _zz__7_27_inner_macOut_2);
  assign _zz__7_27_inner_macOut_2 = (($signed(_zz__7_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_27_inner_activation;
    end else begin
      io_macOut = _7_27_inner_macOut;
    end
  end

  assign _zz__7_27_inner_macOut = ($signed(_zz__zz__7_27_inner_macOut) + $signed(_zz__zz__7_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_27_inner_activation <= 8'h00;
      _7_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_27_inner_activation <= io_addInput;
      end else begin
        _7_27_inner_macOut <= _zz__7_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_250 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_26_inner_macOut;
  wire       [15:0]   _zz__zz__7_26_inner_macOut_1;
  wire       [15:0]   _zz__7_26_inner_macOut_1;
  wire       [15:0]   _zz__7_26_inner_macOut_2;
  reg        [7:0]    _7_26_inner_activation;
  reg        [7:0]    _7_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_26_inner_macOut;

  assign _zz__zz__7_26_inner_macOut = ($signed(io_mulInput) * $signed(_7_26_inner_activation));
  assign _zz__zz__7_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_26_inner_macOut)) ? 16'h007f : _zz__7_26_inner_macOut_2);
  assign _zz__7_26_inner_macOut_2 = (($signed(_zz__7_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_26_inner_activation;
    end else begin
      io_macOut = _7_26_inner_macOut;
    end
  end

  assign _zz__7_26_inner_macOut = ($signed(_zz__zz__7_26_inner_macOut) + $signed(_zz__zz__7_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_26_inner_activation <= 8'h00;
      _7_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_26_inner_activation <= io_addInput;
      end else begin
        _7_26_inner_macOut <= _zz__7_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_249 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_25_inner_macOut;
  wire       [15:0]   _zz__zz__7_25_inner_macOut_1;
  wire       [15:0]   _zz__7_25_inner_macOut_1;
  wire       [15:0]   _zz__7_25_inner_macOut_2;
  reg        [7:0]    _7_25_inner_activation;
  reg        [7:0]    _7_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_25_inner_macOut;

  assign _zz__zz__7_25_inner_macOut = ($signed(io_mulInput) * $signed(_7_25_inner_activation));
  assign _zz__zz__7_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_25_inner_macOut)) ? 16'h007f : _zz__7_25_inner_macOut_2);
  assign _zz__7_25_inner_macOut_2 = (($signed(_zz__7_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_25_inner_activation;
    end else begin
      io_macOut = _7_25_inner_macOut;
    end
  end

  assign _zz__7_25_inner_macOut = ($signed(_zz__zz__7_25_inner_macOut) + $signed(_zz__zz__7_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_25_inner_activation <= 8'h00;
      _7_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_25_inner_activation <= io_addInput;
      end else begin
        _7_25_inner_macOut <= _zz__7_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_248 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_24_inner_macOut;
  wire       [15:0]   _zz__zz__7_24_inner_macOut_1;
  wire       [15:0]   _zz__7_24_inner_macOut_1;
  wire       [15:0]   _zz__7_24_inner_macOut_2;
  reg        [7:0]    _7_24_inner_activation;
  reg        [7:0]    _7_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_24_inner_macOut;

  assign _zz__zz__7_24_inner_macOut = ($signed(io_mulInput) * $signed(_7_24_inner_activation));
  assign _zz__zz__7_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_24_inner_macOut)) ? 16'h007f : _zz__7_24_inner_macOut_2);
  assign _zz__7_24_inner_macOut_2 = (($signed(_zz__7_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_24_inner_activation;
    end else begin
      io_macOut = _7_24_inner_macOut;
    end
  end

  assign _zz__7_24_inner_macOut = ($signed(_zz__zz__7_24_inner_macOut) + $signed(_zz__zz__7_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_24_inner_activation <= 8'h00;
      _7_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_24_inner_activation <= io_addInput;
      end else begin
        _7_24_inner_macOut <= _zz__7_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_247 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_23_inner_macOut;
  wire       [15:0]   _zz__zz__7_23_inner_macOut_1;
  wire       [15:0]   _zz__7_23_inner_macOut_1;
  wire       [15:0]   _zz__7_23_inner_macOut_2;
  reg        [7:0]    _7_23_inner_activation;
  reg        [7:0]    _7_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_23_inner_macOut;

  assign _zz__zz__7_23_inner_macOut = ($signed(io_mulInput) * $signed(_7_23_inner_activation));
  assign _zz__zz__7_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_23_inner_macOut)) ? 16'h007f : _zz__7_23_inner_macOut_2);
  assign _zz__7_23_inner_macOut_2 = (($signed(_zz__7_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_23_inner_activation;
    end else begin
      io_macOut = _7_23_inner_macOut;
    end
  end

  assign _zz__7_23_inner_macOut = ($signed(_zz__zz__7_23_inner_macOut) + $signed(_zz__zz__7_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_23_inner_activation <= 8'h00;
      _7_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_23_inner_activation <= io_addInput;
      end else begin
        _7_23_inner_macOut <= _zz__7_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_246 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_22_inner_macOut;
  wire       [15:0]   _zz__zz__7_22_inner_macOut_1;
  wire       [15:0]   _zz__7_22_inner_macOut_1;
  wire       [15:0]   _zz__7_22_inner_macOut_2;
  reg        [7:0]    _7_22_inner_activation;
  reg        [7:0]    _7_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_22_inner_macOut;

  assign _zz__zz__7_22_inner_macOut = ($signed(io_mulInput) * $signed(_7_22_inner_activation));
  assign _zz__zz__7_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_22_inner_macOut)) ? 16'h007f : _zz__7_22_inner_macOut_2);
  assign _zz__7_22_inner_macOut_2 = (($signed(_zz__7_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_22_inner_activation;
    end else begin
      io_macOut = _7_22_inner_macOut;
    end
  end

  assign _zz__7_22_inner_macOut = ($signed(_zz__zz__7_22_inner_macOut) + $signed(_zz__zz__7_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_22_inner_activation <= 8'h00;
      _7_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_22_inner_activation <= io_addInput;
      end else begin
        _7_22_inner_macOut <= _zz__7_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_245 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_21_inner_macOut;
  wire       [15:0]   _zz__zz__7_21_inner_macOut_1;
  wire       [15:0]   _zz__7_21_inner_macOut_1;
  wire       [15:0]   _zz__7_21_inner_macOut_2;
  reg        [7:0]    _7_21_inner_activation;
  reg        [7:0]    _7_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_21_inner_macOut;

  assign _zz__zz__7_21_inner_macOut = ($signed(io_mulInput) * $signed(_7_21_inner_activation));
  assign _zz__zz__7_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_21_inner_macOut)) ? 16'h007f : _zz__7_21_inner_macOut_2);
  assign _zz__7_21_inner_macOut_2 = (($signed(_zz__7_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_21_inner_activation;
    end else begin
      io_macOut = _7_21_inner_macOut;
    end
  end

  assign _zz__7_21_inner_macOut = ($signed(_zz__zz__7_21_inner_macOut) + $signed(_zz__zz__7_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_21_inner_activation <= 8'h00;
      _7_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_21_inner_activation <= io_addInput;
      end else begin
        _7_21_inner_macOut <= _zz__7_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_244 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_20_inner_macOut;
  wire       [15:0]   _zz__zz__7_20_inner_macOut_1;
  wire       [15:0]   _zz__7_20_inner_macOut_1;
  wire       [15:0]   _zz__7_20_inner_macOut_2;
  reg        [7:0]    _7_20_inner_activation;
  reg        [7:0]    _7_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_20_inner_macOut;

  assign _zz__zz__7_20_inner_macOut = ($signed(io_mulInput) * $signed(_7_20_inner_activation));
  assign _zz__zz__7_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_20_inner_macOut)) ? 16'h007f : _zz__7_20_inner_macOut_2);
  assign _zz__7_20_inner_macOut_2 = (($signed(_zz__7_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_20_inner_activation;
    end else begin
      io_macOut = _7_20_inner_macOut;
    end
  end

  assign _zz__7_20_inner_macOut = ($signed(_zz__zz__7_20_inner_macOut) + $signed(_zz__zz__7_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_20_inner_activation <= 8'h00;
      _7_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_20_inner_activation <= io_addInput;
      end else begin
        _7_20_inner_macOut <= _zz__7_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_243 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_19_inner_macOut;
  wire       [15:0]   _zz__zz__7_19_inner_macOut_1;
  wire       [15:0]   _zz__7_19_inner_macOut_1;
  wire       [15:0]   _zz__7_19_inner_macOut_2;
  reg        [7:0]    _7_19_inner_activation;
  reg        [7:0]    _7_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_19_inner_macOut;

  assign _zz__zz__7_19_inner_macOut = ($signed(io_mulInput) * $signed(_7_19_inner_activation));
  assign _zz__zz__7_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_19_inner_macOut)) ? 16'h007f : _zz__7_19_inner_macOut_2);
  assign _zz__7_19_inner_macOut_2 = (($signed(_zz__7_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_19_inner_activation;
    end else begin
      io_macOut = _7_19_inner_macOut;
    end
  end

  assign _zz__7_19_inner_macOut = ($signed(_zz__zz__7_19_inner_macOut) + $signed(_zz__zz__7_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_19_inner_activation <= 8'h00;
      _7_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_19_inner_activation <= io_addInput;
      end else begin
        _7_19_inner_macOut <= _zz__7_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_242 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_18_inner_macOut;
  wire       [15:0]   _zz__zz__7_18_inner_macOut_1;
  wire       [15:0]   _zz__7_18_inner_macOut_1;
  wire       [15:0]   _zz__7_18_inner_macOut_2;
  reg        [7:0]    _7_18_inner_activation;
  reg        [7:0]    _7_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_18_inner_macOut;

  assign _zz__zz__7_18_inner_macOut = ($signed(io_mulInput) * $signed(_7_18_inner_activation));
  assign _zz__zz__7_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_18_inner_macOut)) ? 16'h007f : _zz__7_18_inner_macOut_2);
  assign _zz__7_18_inner_macOut_2 = (($signed(_zz__7_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_18_inner_activation;
    end else begin
      io_macOut = _7_18_inner_macOut;
    end
  end

  assign _zz__7_18_inner_macOut = ($signed(_zz__zz__7_18_inner_macOut) + $signed(_zz__zz__7_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_18_inner_activation <= 8'h00;
      _7_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_18_inner_activation <= io_addInput;
      end else begin
        _7_18_inner_macOut <= _zz__7_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_241 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_17_inner_macOut;
  wire       [15:0]   _zz__zz__7_17_inner_macOut_1;
  wire       [15:0]   _zz__7_17_inner_macOut_1;
  wire       [15:0]   _zz__7_17_inner_macOut_2;
  reg        [7:0]    _7_17_inner_activation;
  reg        [7:0]    _7_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_17_inner_macOut;

  assign _zz__zz__7_17_inner_macOut = ($signed(io_mulInput) * $signed(_7_17_inner_activation));
  assign _zz__zz__7_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_17_inner_macOut)) ? 16'h007f : _zz__7_17_inner_macOut_2);
  assign _zz__7_17_inner_macOut_2 = (($signed(_zz__7_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_17_inner_activation;
    end else begin
      io_macOut = _7_17_inner_macOut;
    end
  end

  assign _zz__7_17_inner_macOut = ($signed(_zz__zz__7_17_inner_macOut) + $signed(_zz__zz__7_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_17_inner_activation <= 8'h00;
      _7_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_17_inner_activation <= io_addInput;
      end else begin
        _7_17_inner_macOut <= _zz__7_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_240 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_16_inner_macOut;
  wire       [15:0]   _zz__zz__7_16_inner_macOut_1;
  wire       [15:0]   _zz__7_16_inner_macOut_1;
  wire       [15:0]   _zz__7_16_inner_macOut_2;
  reg        [7:0]    _7_16_inner_activation;
  reg        [7:0]    _7_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_16_inner_macOut;

  assign _zz__zz__7_16_inner_macOut = ($signed(io_mulInput) * $signed(_7_16_inner_activation));
  assign _zz__zz__7_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_16_inner_macOut)) ? 16'h007f : _zz__7_16_inner_macOut_2);
  assign _zz__7_16_inner_macOut_2 = (($signed(_zz__7_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_16_inner_activation;
    end else begin
      io_macOut = _7_16_inner_macOut;
    end
  end

  assign _zz__7_16_inner_macOut = ($signed(_zz__zz__7_16_inner_macOut) + $signed(_zz__zz__7_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_16_inner_activation <= 8'h00;
      _7_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_16_inner_activation <= io_addInput;
      end else begin
        _7_16_inner_macOut <= _zz__7_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_239 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_15_inner_macOut;
  wire       [15:0]   _zz__zz__7_15_inner_macOut_1;
  wire       [15:0]   _zz__7_15_inner_macOut_1;
  wire       [15:0]   _zz__7_15_inner_macOut_2;
  reg        [7:0]    _7_15_inner_activation;
  reg        [7:0]    _7_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_15_inner_macOut;

  assign _zz__zz__7_15_inner_macOut = ($signed(io_mulInput) * $signed(_7_15_inner_activation));
  assign _zz__zz__7_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_15_inner_macOut)) ? 16'h007f : _zz__7_15_inner_macOut_2);
  assign _zz__7_15_inner_macOut_2 = (($signed(_zz__7_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_15_inner_activation;
    end else begin
      io_macOut = _7_15_inner_macOut;
    end
  end

  assign _zz__7_15_inner_macOut = ($signed(_zz__zz__7_15_inner_macOut) + $signed(_zz__zz__7_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_15_inner_activation <= 8'h00;
      _7_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_15_inner_activation <= io_addInput;
      end else begin
        _7_15_inner_macOut <= _zz__7_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_238 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_14_inner_macOut;
  wire       [15:0]   _zz__zz__7_14_inner_macOut_1;
  wire       [15:0]   _zz__7_14_inner_macOut_1;
  wire       [15:0]   _zz__7_14_inner_macOut_2;
  reg        [7:0]    _7_14_inner_activation;
  reg        [7:0]    _7_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_14_inner_macOut;

  assign _zz__zz__7_14_inner_macOut = ($signed(io_mulInput) * $signed(_7_14_inner_activation));
  assign _zz__zz__7_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_14_inner_macOut)) ? 16'h007f : _zz__7_14_inner_macOut_2);
  assign _zz__7_14_inner_macOut_2 = (($signed(_zz__7_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_14_inner_activation;
    end else begin
      io_macOut = _7_14_inner_macOut;
    end
  end

  assign _zz__7_14_inner_macOut = ($signed(_zz__zz__7_14_inner_macOut) + $signed(_zz__zz__7_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_14_inner_activation <= 8'h00;
      _7_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_14_inner_activation <= io_addInput;
      end else begin
        _7_14_inner_macOut <= _zz__7_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_237 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_13_inner_macOut;
  wire       [15:0]   _zz__zz__7_13_inner_macOut_1;
  wire       [15:0]   _zz__7_13_inner_macOut_1;
  wire       [15:0]   _zz__7_13_inner_macOut_2;
  reg        [7:0]    _7_13_inner_activation;
  reg        [7:0]    _7_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_13_inner_macOut;

  assign _zz__zz__7_13_inner_macOut = ($signed(io_mulInput) * $signed(_7_13_inner_activation));
  assign _zz__zz__7_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_13_inner_macOut)) ? 16'h007f : _zz__7_13_inner_macOut_2);
  assign _zz__7_13_inner_macOut_2 = (($signed(_zz__7_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_13_inner_activation;
    end else begin
      io_macOut = _7_13_inner_macOut;
    end
  end

  assign _zz__7_13_inner_macOut = ($signed(_zz__zz__7_13_inner_macOut) + $signed(_zz__zz__7_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_13_inner_activation <= 8'h00;
      _7_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_13_inner_activation <= io_addInput;
      end else begin
        _7_13_inner_macOut <= _zz__7_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_236 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_12_inner_macOut;
  wire       [15:0]   _zz__zz__7_12_inner_macOut_1;
  wire       [15:0]   _zz__7_12_inner_macOut_1;
  wire       [15:0]   _zz__7_12_inner_macOut_2;
  reg        [7:0]    _7_12_inner_activation;
  reg        [7:0]    _7_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_12_inner_macOut;

  assign _zz__zz__7_12_inner_macOut = ($signed(io_mulInput) * $signed(_7_12_inner_activation));
  assign _zz__zz__7_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_12_inner_macOut)) ? 16'h007f : _zz__7_12_inner_macOut_2);
  assign _zz__7_12_inner_macOut_2 = (($signed(_zz__7_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_12_inner_activation;
    end else begin
      io_macOut = _7_12_inner_macOut;
    end
  end

  assign _zz__7_12_inner_macOut = ($signed(_zz__zz__7_12_inner_macOut) + $signed(_zz__zz__7_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_12_inner_activation <= 8'h00;
      _7_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_12_inner_activation <= io_addInput;
      end else begin
        _7_12_inner_macOut <= _zz__7_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_235 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_11_inner_macOut;
  wire       [15:0]   _zz__zz__7_11_inner_macOut_1;
  wire       [15:0]   _zz__7_11_inner_macOut_1;
  wire       [15:0]   _zz__7_11_inner_macOut_2;
  reg        [7:0]    _7_11_inner_activation;
  reg        [7:0]    _7_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_11_inner_macOut;

  assign _zz__zz__7_11_inner_macOut = ($signed(io_mulInput) * $signed(_7_11_inner_activation));
  assign _zz__zz__7_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_11_inner_macOut)) ? 16'h007f : _zz__7_11_inner_macOut_2);
  assign _zz__7_11_inner_macOut_2 = (($signed(_zz__7_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_11_inner_activation;
    end else begin
      io_macOut = _7_11_inner_macOut;
    end
  end

  assign _zz__7_11_inner_macOut = ($signed(_zz__zz__7_11_inner_macOut) + $signed(_zz__zz__7_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_11_inner_activation <= 8'h00;
      _7_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_11_inner_activation <= io_addInput;
      end else begin
        _7_11_inner_macOut <= _zz__7_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_234 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_10_inner_macOut;
  wire       [15:0]   _zz__zz__7_10_inner_macOut_1;
  wire       [15:0]   _zz__7_10_inner_macOut_1;
  wire       [15:0]   _zz__7_10_inner_macOut_2;
  reg        [7:0]    _7_10_inner_activation;
  reg        [7:0]    _7_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_10_inner_macOut;

  assign _zz__zz__7_10_inner_macOut = ($signed(io_mulInput) * $signed(_7_10_inner_activation));
  assign _zz__zz__7_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_10_inner_macOut)) ? 16'h007f : _zz__7_10_inner_macOut_2);
  assign _zz__7_10_inner_macOut_2 = (($signed(_zz__7_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_10_inner_activation;
    end else begin
      io_macOut = _7_10_inner_macOut;
    end
  end

  assign _zz__7_10_inner_macOut = ($signed(_zz__zz__7_10_inner_macOut) + $signed(_zz__zz__7_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_10_inner_activation <= 8'h00;
      _7_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_10_inner_activation <= io_addInput;
      end else begin
        _7_10_inner_macOut <= _zz__7_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_233 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_9_inner_macOut;
  wire       [15:0]   _zz__zz__7_9_inner_macOut_1;
  wire       [15:0]   _zz__7_9_inner_macOut_1;
  wire       [15:0]   _zz__7_9_inner_macOut_2;
  reg        [7:0]    _7_9_inner_activation;
  reg        [7:0]    _7_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_9_inner_macOut;

  assign _zz__zz__7_9_inner_macOut = ($signed(io_mulInput) * $signed(_7_9_inner_activation));
  assign _zz__zz__7_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_9_inner_macOut)) ? 16'h007f : _zz__7_9_inner_macOut_2);
  assign _zz__7_9_inner_macOut_2 = (($signed(_zz__7_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_9_inner_activation;
    end else begin
      io_macOut = _7_9_inner_macOut;
    end
  end

  assign _zz__7_9_inner_macOut = ($signed(_zz__zz__7_9_inner_macOut) + $signed(_zz__zz__7_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_9_inner_activation <= 8'h00;
      _7_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_9_inner_activation <= io_addInput;
      end else begin
        _7_9_inner_macOut <= _zz__7_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_232 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_8_inner_macOut;
  wire       [15:0]   _zz__zz__7_8_inner_macOut_1;
  wire       [15:0]   _zz__7_8_inner_macOut_1;
  wire       [15:0]   _zz__7_8_inner_macOut_2;
  reg        [7:0]    _7_8_inner_activation;
  reg        [7:0]    _7_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_8_inner_macOut;

  assign _zz__zz__7_8_inner_macOut = ($signed(io_mulInput) * $signed(_7_8_inner_activation));
  assign _zz__zz__7_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_8_inner_macOut)) ? 16'h007f : _zz__7_8_inner_macOut_2);
  assign _zz__7_8_inner_macOut_2 = (($signed(_zz__7_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_8_inner_activation;
    end else begin
      io_macOut = _7_8_inner_macOut;
    end
  end

  assign _zz__7_8_inner_macOut = ($signed(_zz__zz__7_8_inner_macOut) + $signed(_zz__zz__7_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_8_inner_activation <= 8'h00;
      _7_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_8_inner_activation <= io_addInput;
      end else begin
        _7_8_inner_macOut <= _zz__7_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_231 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_7_inner_macOut;
  wire       [15:0]   _zz__zz__7_7_inner_macOut_1;
  wire       [15:0]   _zz__7_7_inner_macOut_1;
  wire       [15:0]   _zz__7_7_inner_macOut_2;
  reg        [7:0]    _7_7_inner_activation;
  reg        [7:0]    _7_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_7_inner_macOut;

  assign _zz__zz__7_7_inner_macOut = ($signed(io_mulInput) * $signed(_7_7_inner_activation));
  assign _zz__zz__7_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_7_inner_macOut)) ? 16'h007f : _zz__7_7_inner_macOut_2);
  assign _zz__7_7_inner_macOut_2 = (($signed(_zz__7_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_7_inner_activation;
    end else begin
      io_macOut = _7_7_inner_macOut;
    end
  end

  assign _zz__7_7_inner_macOut = ($signed(_zz__zz__7_7_inner_macOut) + $signed(_zz__zz__7_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_7_inner_activation <= 8'h00;
      _7_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_7_inner_activation <= io_addInput;
      end else begin
        _7_7_inner_macOut <= _zz__7_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_230 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_6_inner_macOut;
  wire       [15:0]   _zz__zz__7_6_inner_macOut_1;
  wire       [15:0]   _zz__7_6_inner_macOut_1;
  wire       [15:0]   _zz__7_6_inner_macOut_2;
  reg        [7:0]    _7_6_inner_activation;
  reg        [7:0]    _7_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_6_inner_macOut;

  assign _zz__zz__7_6_inner_macOut = ($signed(io_mulInput) * $signed(_7_6_inner_activation));
  assign _zz__zz__7_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_6_inner_macOut)) ? 16'h007f : _zz__7_6_inner_macOut_2);
  assign _zz__7_6_inner_macOut_2 = (($signed(_zz__7_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_6_inner_activation;
    end else begin
      io_macOut = _7_6_inner_macOut;
    end
  end

  assign _zz__7_6_inner_macOut = ($signed(_zz__zz__7_6_inner_macOut) + $signed(_zz__zz__7_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_6_inner_activation <= 8'h00;
      _7_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_6_inner_activation <= io_addInput;
      end else begin
        _7_6_inner_macOut <= _zz__7_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_229 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_5_inner_macOut;
  wire       [15:0]   _zz__zz__7_5_inner_macOut_1;
  wire       [15:0]   _zz__7_5_inner_macOut_1;
  wire       [15:0]   _zz__7_5_inner_macOut_2;
  reg        [7:0]    _7_5_inner_activation;
  reg        [7:0]    _7_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_5_inner_macOut;

  assign _zz__zz__7_5_inner_macOut = ($signed(io_mulInput) * $signed(_7_5_inner_activation));
  assign _zz__zz__7_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_5_inner_macOut)) ? 16'h007f : _zz__7_5_inner_macOut_2);
  assign _zz__7_5_inner_macOut_2 = (($signed(_zz__7_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_5_inner_activation;
    end else begin
      io_macOut = _7_5_inner_macOut;
    end
  end

  assign _zz__7_5_inner_macOut = ($signed(_zz__zz__7_5_inner_macOut) + $signed(_zz__zz__7_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_5_inner_activation <= 8'h00;
      _7_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_5_inner_activation <= io_addInput;
      end else begin
        _7_5_inner_macOut <= _zz__7_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_228 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_4_inner_macOut;
  wire       [15:0]   _zz__zz__7_4_inner_macOut_1;
  wire       [15:0]   _zz__7_4_inner_macOut_1;
  wire       [15:0]   _zz__7_4_inner_macOut_2;
  reg        [7:0]    _7_4_inner_activation;
  reg        [7:0]    _7_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_4_inner_macOut;

  assign _zz__zz__7_4_inner_macOut = ($signed(io_mulInput) * $signed(_7_4_inner_activation));
  assign _zz__zz__7_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_4_inner_macOut)) ? 16'h007f : _zz__7_4_inner_macOut_2);
  assign _zz__7_4_inner_macOut_2 = (($signed(_zz__7_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_4_inner_activation;
    end else begin
      io_macOut = _7_4_inner_macOut;
    end
  end

  assign _zz__7_4_inner_macOut = ($signed(_zz__zz__7_4_inner_macOut) + $signed(_zz__zz__7_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_4_inner_activation <= 8'h00;
      _7_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_4_inner_activation <= io_addInput;
      end else begin
        _7_4_inner_macOut <= _zz__7_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_227 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_3_inner_macOut;
  wire       [15:0]   _zz__zz__7_3_inner_macOut_1;
  wire       [15:0]   _zz__7_3_inner_macOut_1;
  wire       [15:0]   _zz__7_3_inner_macOut_2;
  reg        [7:0]    _7_3_inner_activation;
  reg        [7:0]    _7_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_3_inner_macOut;

  assign _zz__zz__7_3_inner_macOut = ($signed(io_mulInput) * $signed(_7_3_inner_activation));
  assign _zz__zz__7_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_3_inner_macOut)) ? 16'h007f : _zz__7_3_inner_macOut_2);
  assign _zz__7_3_inner_macOut_2 = (($signed(_zz__7_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_3_inner_activation;
    end else begin
      io_macOut = _7_3_inner_macOut;
    end
  end

  assign _zz__7_3_inner_macOut = ($signed(_zz__zz__7_3_inner_macOut) + $signed(_zz__zz__7_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_3_inner_activation <= 8'h00;
      _7_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_3_inner_activation <= io_addInput;
      end else begin
        _7_3_inner_macOut <= _zz__7_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_226 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_2_inner_macOut;
  wire       [15:0]   _zz__zz__7_2_inner_macOut_1;
  wire       [15:0]   _zz__7_2_inner_macOut_1;
  wire       [15:0]   _zz__7_2_inner_macOut_2;
  reg        [7:0]    _7_2_inner_activation;
  reg        [7:0]    _7_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_2_inner_macOut;

  assign _zz__zz__7_2_inner_macOut = ($signed(io_mulInput) * $signed(_7_2_inner_activation));
  assign _zz__zz__7_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_2_inner_macOut)) ? 16'h007f : _zz__7_2_inner_macOut_2);
  assign _zz__7_2_inner_macOut_2 = (($signed(_zz__7_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_2_inner_activation;
    end else begin
      io_macOut = _7_2_inner_macOut;
    end
  end

  assign _zz__7_2_inner_macOut = ($signed(_zz__zz__7_2_inner_macOut) + $signed(_zz__zz__7_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_2_inner_activation <= 8'h00;
      _7_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_2_inner_activation <= io_addInput;
      end else begin
        _7_2_inner_macOut <= _zz__7_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_225 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_1_inner_macOut;
  wire       [15:0]   _zz__zz__7_1_inner_macOut_1;
  wire       [15:0]   _zz__7_1_inner_macOut_1;
  wire       [15:0]   _zz__7_1_inner_macOut_2;
  reg        [7:0]    _7_1_inner_activation;
  reg        [7:0]    _7_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_1_inner_macOut;

  assign _zz__zz__7_1_inner_macOut = ($signed(io_mulInput) * $signed(_7_1_inner_activation));
  assign _zz__zz__7_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_1_inner_macOut)) ? 16'h007f : _zz__7_1_inner_macOut_2);
  assign _zz__7_1_inner_macOut_2 = (($signed(_zz__7_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_1_inner_activation;
    end else begin
      io_macOut = _7_1_inner_macOut;
    end
  end

  assign _zz__7_1_inner_macOut = ($signed(_zz__zz__7_1_inner_macOut) + $signed(_zz__zz__7_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_1_inner_activation <= 8'h00;
      _7_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_1_inner_activation <= io_addInput;
      end else begin
        _7_1_inner_macOut <= _zz__7_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_224 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__7_0_inner_macOut;
  wire       [15:0]   _zz__zz__7_0_inner_macOut_1;
  wire       [15:0]   _zz__7_0_inner_macOut_1;
  wire       [15:0]   _zz__7_0_inner_macOut_2;
  reg        [7:0]    _7_0_inner_activation;
  reg        [7:0]    _7_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__7_0_inner_macOut;

  assign _zz__zz__7_0_inner_macOut = ($signed(io_mulInput) * $signed(_7_0_inner_activation));
  assign _zz__zz__7_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__7_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__7_0_inner_macOut)) ? 16'h007f : _zz__7_0_inner_macOut_2);
  assign _zz__7_0_inner_macOut_2 = (($signed(_zz__7_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__7_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _7_0_inner_activation;
    end else begin
      io_macOut = _7_0_inner_macOut;
    end
  end

  assign _zz__7_0_inner_macOut = ($signed(_zz__zz__7_0_inner_macOut) + $signed(_zz__zz__7_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _7_0_inner_activation <= 8'h00;
      _7_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _7_0_inner_activation <= io_addInput;
      end else begin
        _7_0_inner_macOut <= _zz__7_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_223 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_31_inner_macOut;
  wire       [15:0]   _zz__zz__6_31_inner_macOut_1;
  wire       [15:0]   _zz__6_31_inner_macOut_1;
  wire       [15:0]   _zz__6_31_inner_macOut_2;
  reg        [7:0]    _6_31_inner_activation;
  reg        [7:0]    _6_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_31_inner_macOut;

  assign _zz__zz__6_31_inner_macOut = ($signed(io_mulInput) * $signed(_6_31_inner_activation));
  assign _zz__zz__6_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_31_inner_macOut)) ? 16'h007f : _zz__6_31_inner_macOut_2);
  assign _zz__6_31_inner_macOut_2 = (($signed(_zz__6_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_31_inner_activation;
    end else begin
      io_macOut = _6_31_inner_macOut;
    end
  end

  assign _zz__6_31_inner_macOut = ($signed(_zz__zz__6_31_inner_macOut) + $signed(_zz__zz__6_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_31_inner_activation <= 8'h00;
      _6_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_31_inner_activation <= io_addInput;
      end else begin
        _6_31_inner_macOut <= _zz__6_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_222 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_30_inner_macOut;
  wire       [15:0]   _zz__zz__6_30_inner_macOut_1;
  wire       [15:0]   _zz__6_30_inner_macOut_1;
  wire       [15:0]   _zz__6_30_inner_macOut_2;
  reg        [7:0]    _6_30_inner_activation;
  reg        [7:0]    _6_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_30_inner_macOut;

  assign _zz__zz__6_30_inner_macOut = ($signed(io_mulInput) * $signed(_6_30_inner_activation));
  assign _zz__zz__6_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_30_inner_macOut)) ? 16'h007f : _zz__6_30_inner_macOut_2);
  assign _zz__6_30_inner_macOut_2 = (($signed(_zz__6_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_30_inner_activation;
    end else begin
      io_macOut = _6_30_inner_macOut;
    end
  end

  assign _zz__6_30_inner_macOut = ($signed(_zz__zz__6_30_inner_macOut) + $signed(_zz__zz__6_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_30_inner_activation <= 8'h00;
      _6_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_30_inner_activation <= io_addInput;
      end else begin
        _6_30_inner_macOut <= _zz__6_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_221 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_29_inner_macOut;
  wire       [15:0]   _zz__zz__6_29_inner_macOut_1;
  wire       [15:0]   _zz__6_29_inner_macOut_1;
  wire       [15:0]   _zz__6_29_inner_macOut_2;
  reg        [7:0]    _6_29_inner_activation;
  reg        [7:0]    _6_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_29_inner_macOut;

  assign _zz__zz__6_29_inner_macOut = ($signed(io_mulInput) * $signed(_6_29_inner_activation));
  assign _zz__zz__6_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_29_inner_macOut)) ? 16'h007f : _zz__6_29_inner_macOut_2);
  assign _zz__6_29_inner_macOut_2 = (($signed(_zz__6_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_29_inner_activation;
    end else begin
      io_macOut = _6_29_inner_macOut;
    end
  end

  assign _zz__6_29_inner_macOut = ($signed(_zz__zz__6_29_inner_macOut) + $signed(_zz__zz__6_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_29_inner_activation <= 8'h00;
      _6_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_29_inner_activation <= io_addInput;
      end else begin
        _6_29_inner_macOut <= _zz__6_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_220 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_28_inner_macOut;
  wire       [15:0]   _zz__zz__6_28_inner_macOut_1;
  wire       [15:0]   _zz__6_28_inner_macOut_1;
  wire       [15:0]   _zz__6_28_inner_macOut_2;
  reg        [7:0]    _6_28_inner_activation;
  reg        [7:0]    _6_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_28_inner_macOut;

  assign _zz__zz__6_28_inner_macOut = ($signed(io_mulInput) * $signed(_6_28_inner_activation));
  assign _zz__zz__6_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_28_inner_macOut)) ? 16'h007f : _zz__6_28_inner_macOut_2);
  assign _zz__6_28_inner_macOut_2 = (($signed(_zz__6_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_28_inner_activation;
    end else begin
      io_macOut = _6_28_inner_macOut;
    end
  end

  assign _zz__6_28_inner_macOut = ($signed(_zz__zz__6_28_inner_macOut) + $signed(_zz__zz__6_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_28_inner_activation <= 8'h00;
      _6_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_28_inner_activation <= io_addInput;
      end else begin
        _6_28_inner_macOut <= _zz__6_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_219 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_27_inner_macOut;
  wire       [15:0]   _zz__zz__6_27_inner_macOut_1;
  wire       [15:0]   _zz__6_27_inner_macOut_1;
  wire       [15:0]   _zz__6_27_inner_macOut_2;
  reg        [7:0]    _6_27_inner_activation;
  reg        [7:0]    _6_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_27_inner_macOut;

  assign _zz__zz__6_27_inner_macOut = ($signed(io_mulInput) * $signed(_6_27_inner_activation));
  assign _zz__zz__6_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_27_inner_macOut)) ? 16'h007f : _zz__6_27_inner_macOut_2);
  assign _zz__6_27_inner_macOut_2 = (($signed(_zz__6_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_27_inner_activation;
    end else begin
      io_macOut = _6_27_inner_macOut;
    end
  end

  assign _zz__6_27_inner_macOut = ($signed(_zz__zz__6_27_inner_macOut) + $signed(_zz__zz__6_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_27_inner_activation <= 8'h00;
      _6_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_27_inner_activation <= io_addInput;
      end else begin
        _6_27_inner_macOut <= _zz__6_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_218 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_26_inner_macOut;
  wire       [15:0]   _zz__zz__6_26_inner_macOut_1;
  wire       [15:0]   _zz__6_26_inner_macOut_1;
  wire       [15:0]   _zz__6_26_inner_macOut_2;
  reg        [7:0]    _6_26_inner_activation;
  reg        [7:0]    _6_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_26_inner_macOut;

  assign _zz__zz__6_26_inner_macOut = ($signed(io_mulInput) * $signed(_6_26_inner_activation));
  assign _zz__zz__6_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_26_inner_macOut)) ? 16'h007f : _zz__6_26_inner_macOut_2);
  assign _zz__6_26_inner_macOut_2 = (($signed(_zz__6_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_26_inner_activation;
    end else begin
      io_macOut = _6_26_inner_macOut;
    end
  end

  assign _zz__6_26_inner_macOut = ($signed(_zz__zz__6_26_inner_macOut) + $signed(_zz__zz__6_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_26_inner_activation <= 8'h00;
      _6_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_26_inner_activation <= io_addInput;
      end else begin
        _6_26_inner_macOut <= _zz__6_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_217 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_25_inner_macOut;
  wire       [15:0]   _zz__zz__6_25_inner_macOut_1;
  wire       [15:0]   _zz__6_25_inner_macOut_1;
  wire       [15:0]   _zz__6_25_inner_macOut_2;
  reg        [7:0]    _6_25_inner_activation;
  reg        [7:0]    _6_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_25_inner_macOut;

  assign _zz__zz__6_25_inner_macOut = ($signed(io_mulInput) * $signed(_6_25_inner_activation));
  assign _zz__zz__6_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_25_inner_macOut)) ? 16'h007f : _zz__6_25_inner_macOut_2);
  assign _zz__6_25_inner_macOut_2 = (($signed(_zz__6_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_25_inner_activation;
    end else begin
      io_macOut = _6_25_inner_macOut;
    end
  end

  assign _zz__6_25_inner_macOut = ($signed(_zz__zz__6_25_inner_macOut) + $signed(_zz__zz__6_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_25_inner_activation <= 8'h00;
      _6_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_25_inner_activation <= io_addInput;
      end else begin
        _6_25_inner_macOut <= _zz__6_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_216 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_24_inner_macOut;
  wire       [15:0]   _zz__zz__6_24_inner_macOut_1;
  wire       [15:0]   _zz__6_24_inner_macOut_1;
  wire       [15:0]   _zz__6_24_inner_macOut_2;
  reg        [7:0]    _6_24_inner_activation;
  reg        [7:0]    _6_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_24_inner_macOut;

  assign _zz__zz__6_24_inner_macOut = ($signed(io_mulInput) * $signed(_6_24_inner_activation));
  assign _zz__zz__6_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_24_inner_macOut)) ? 16'h007f : _zz__6_24_inner_macOut_2);
  assign _zz__6_24_inner_macOut_2 = (($signed(_zz__6_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_24_inner_activation;
    end else begin
      io_macOut = _6_24_inner_macOut;
    end
  end

  assign _zz__6_24_inner_macOut = ($signed(_zz__zz__6_24_inner_macOut) + $signed(_zz__zz__6_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_24_inner_activation <= 8'h00;
      _6_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_24_inner_activation <= io_addInput;
      end else begin
        _6_24_inner_macOut <= _zz__6_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_215 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_23_inner_macOut;
  wire       [15:0]   _zz__zz__6_23_inner_macOut_1;
  wire       [15:0]   _zz__6_23_inner_macOut_1;
  wire       [15:0]   _zz__6_23_inner_macOut_2;
  reg        [7:0]    _6_23_inner_activation;
  reg        [7:0]    _6_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_23_inner_macOut;

  assign _zz__zz__6_23_inner_macOut = ($signed(io_mulInput) * $signed(_6_23_inner_activation));
  assign _zz__zz__6_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_23_inner_macOut)) ? 16'h007f : _zz__6_23_inner_macOut_2);
  assign _zz__6_23_inner_macOut_2 = (($signed(_zz__6_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_23_inner_activation;
    end else begin
      io_macOut = _6_23_inner_macOut;
    end
  end

  assign _zz__6_23_inner_macOut = ($signed(_zz__zz__6_23_inner_macOut) + $signed(_zz__zz__6_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_23_inner_activation <= 8'h00;
      _6_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_23_inner_activation <= io_addInput;
      end else begin
        _6_23_inner_macOut <= _zz__6_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_214 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_22_inner_macOut;
  wire       [15:0]   _zz__zz__6_22_inner_macOut_1;
  wire       [15:0]   _zz__6_22_inner_macOut_1;
  wire       [15:0]   _zz__6_22_inner_macOut_2;
  reg        [7:0]    _6_22_inner_activation;
  reg        [7:0]    _6_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_22_inner_macOut;

  assign _zz__zz__6_22_inner_macOut = ($signed(io_mulInput) * $signed(_6_22_inner_activation));
  assign _zz__zz__6_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_22_inner_macOut)) ? 16'h007f : _zz__6_22_inner_macOut_2);
  assign _zz__6_22_inner_macOut_2 = (($signed(_zz__6_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_22_inner_activation;
    end else begin
      io_macOut = _6_22_inner_macOut;
    end
  end

  assign _zz__6_22_inner_macOut = ($signed(_zz__zz__6_22_inner_macOut) + $signed(_zz__zz__6_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_22_inner_activation <= 8'h00;
      _6_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_22_inner_activation <= io_addInput;
      end else begin
        _6_22_inner_macOut <= _zz__6_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_213 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_21_inner_macOut;
  wire       [15:0]   _zz__zz__6_21_inner_macOut_1;
  wire       [15:0]   _zz__6_21_inner_macOut_1;
  wire       [15:0]   _zz__6_21_inner_macOut_2;
  reg        [7:0]    _6_21_inner_activation;
  reg        [7:0]    _6_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_21_inner_macOut;

  assign _zz__zz__6_21_inner_macOut = ($signed(io_mulInput) * $signed(_6_21_inner_activation));
  assign _zz__zz__6_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_21_inner_macOut)) ? 16'h007f : _zz__6_21_inner_macOut_2);
  assign _zz__6_21_inner_macOut_2 = (($signed(_zz__6_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_21_inner_activation;
    end else begin
      io_macOut = _6_21_inner_macOut;
    end
  end

  assign _zz__6_21_inner_macOut = ($signed(_zz__zz__6_21_inner_macOut) + $signed(_zz__zz__6_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_21_inner_activation <= 8'h00;
      _6_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_21_inner_activation <= io_addInput;
      end else begin
        _6_21_inner_macOut <= _zz__6_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_212 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_20_inner_macOut;
  wire       [15:0]   _zz__zz__6_20_inner_macOut_1;
  wire       [15:0]   _zz__6_20_inner_macOut_1;
  wire       [15:0]   _zz__6_20_inner_macOut_2;
  reg        [7:0]    _6_20_inner_activation;
  reg        [7:0]    _6_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_20_inner_macOut;

  assign _zz__zz__6_20_inner_macOut = ($signed(io_mulInput) * $signed(_6_20_inner_activation));
  assign _zz__zz__6_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_20_inner_macOut)) ? 16'h007f : _zz__6_20_inner_macOut_2);
  assign _zz__6_20_inner_macOut_2 = (($signed(_zz__6_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_20_inner_activation;
    end else begin
      io_macOut = _6_20_inner_macOut;
    end
  end

  assign _zz__6_20_inner_macOut = ($signed(_zz__zz__6_20_inner_macOut) + $signed(_zz__zz__6_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_20_inner_activation <= 8'h00;
      _6_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_20_inner_activation <= io_addInput;
      end else begin
        _6_20_inner_macOut <= _zz__6_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_211 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_19_inner_macOut;
  wire       [15:0]   _zz__zz__6_19_inner_macOut_1;
  wire       [15:0]   _zz__6_19_inner_macOut_1;
  wire       [15:0]   _zz__6_19_inner_macOut_2;
  reg        [7:0]    _6_19_inner_activation;
  reg        [7:0]    _6_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_19_inner_macOut;

  assign _zz__zz__6_19_inner_macOut = ($signed(io_mulInput) * $signed(_6_19_inner_activation));
  assign _zz__zz__6_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_19_inner_macOut)) ? 16'h007f : _zz__6_19_inner_macOut_2);
  assign _zz__6_19_inner_macOut_2 = (($signed(_zz__6_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_19_inner_activation;
    end else begin
      io_macOut = _6_19_inner_macOut;
    end
  end

  assign _zz__6_19_inner_macOut = ($signed(_zz__zz__6_19_inner_macOut) + $signed(_zz__zz__6_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_19_inner_activation <= 8'h00;
      _6_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_19_inner_activation <= io_addInput;
      end else begin
        _6_19_inner_macOut <= _zz__6_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_210 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_18_inner_macOut;
  wire       [15:0]   _zz__zz__6_18_inner_macOut_1;
  wire       [15:0]   _zz__6_18_inner_macOut_1;
  wire       [15:0]   _zz__6_18_inner_macOut_2;
  reg        [7:0]    _6_18_inner_activation;
  reg        [7:0]    _6_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_18_inner_macOut;

  assign _zz__zz__6_18_inner_macOut = ($signed(io_mulInput) * $signed(_6_18_inner_activation));
  assign _zz__zz__6_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_18_inner_macOut)) ? 16'h007f : _zz__6_18_inner_macOut_2);
  assign _zz__6_18_inner_macOut_2 = (($signed(_zz__6_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_18_inner_activation;
    end else begin
      io_macOut = _6_18_inner_macOut;
    end
  end

  assign _zz__6_18_inner_macOut = ($signed(_zz__zz__6_18_inner_macOut) + $signed(_zz__zz__6_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_18_inner_activation <= 8'h00;
      _6_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_18_inner_activation <= io_addInput;
      end else begin
        _6_18_inner_macOut <= _zz__6_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_209 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_17_inner_macOut;
  wire       [15:0]   _zz__zz__6_17_inner_macOut_1;
  wire       [15:0]   _zz__6_17_inner_macOut_1;
  wire       [15:0]   _zz__6_17_inner_macOut_2;
  reg        [7:0]    _6_17_inner_activation;
  reg        [7:0]    _6_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_17_inner_macOut;

  assign _zz__zz__6_17_inner_macOut = ($signed(io_mulInput) * $signed(_6_17_inner_activation));
  assign _zz__zz__6_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_17_inner_macOut)) ? 16'h007f : _zz__6_17_inner_macOut_2);
  assign _zz__6_17_inner_macOut_2 = (($signed(_zz__6_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_17_inner_activation;
    end else begin
      io_macOut = _6_17_inner_macOut;
    end
  end

  assign _zz__6_17_inner_macOut = ($signed(_zz__zz__6_17_inner_macOut) + $signed(_zz__zz__6_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_17_inner_activation <= 8'h00;
      _6_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_17_inner_activation <= io_addInput;
      end else begin
        _6_17_inner_macOut <= _zz__6_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_208 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_16_inner_macOut;
  wire       [15:0]   _zz__zz__6_16_inner_macOut_1;
  wire       [15:0]   _zz__6_16_inner_macOut_1;
  wire       [15:0]   _zz__6_16_inner_macOut_2;
  reg        [7:0]    _6_16_inner_activation;
  reg        [7:0]    _6_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_16_inner_macOut;

  assign _zz__zz__6_16_inner_macOut = ($signed(io_mulInput) * $signed(_6_16_inner_activation));
  assign _zz__zz__6_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_16_inner_macOut)) ? 16'h007f : _zz__6_16_inner_macOut_2);
  assign _zz__6_16_inner_macOut_2 = (($signed(_zz__6_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_16_inner_activation;
    end else begin
      io_macOut = _6_16_inner_macOut;
    end
  end

  assign _zz__6_16_inner_macOut = ($signed(_zz__zz__6_16_inner_macOut) + $signed(_zz__zz__6_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_16_inner_activation <= 8'h00;
      _6_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_16_inner_activation <= io_addInput;
      end else begin
        _6_16_inner_macOut <= _zz__6_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_207 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_15_inner_macOut;
  wire       [15:0]   _zz__zz__6_15_inner_macOut_1;
  wire       [15:0]   _zz__6_15_inner_macOut_1;
  wire       [15:0]   _zz__6_15_inner_macOut_2;
  reg        [7:0]    _6_15_inner_activation;
  reg        [7:0]    _6_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_15_inner_macOut;

  assign _zz__zz__6_15_inner_macOut = ($signed(io_mulInput) * $signed(_6_15_inner_activation));
  assign _zz__zz__6_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_15_inner_macOut)) ? 16'h007f : _zz__6_15_inner_macOut_2);
  assign _zz__6_15_inner_macOut_2 = (($signed(_zz__6_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_15_inner_activation;
    end else begin
      io_macOut = _6_15_inner_macOut;
    end
  end

  assign _zz__6_15_inner_macOut = ($signed(_zz__zz__6_15_inner_macOut) + $signed(_zz__zz__6_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_15_inner_activation <= 8'h00;
      _6_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_15_inner_activation <= io_addInput;
      end else begin
        _6_15_inner_macOut <= _zz__6_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_206 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_14_inner_macOut;
  wire       [15:0]   _zz__zz__6_14_inner_macOut_1;
  wire       [15:0]   _zz__6_14_inner_macOut_1;
  wire       [15:0]   _zz__6_14_inner_macOut_2;
  reg        [7:0]    _6_14_inner_activation;
  reg        [7:0]    _6_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_14_inner_macOut;

  assign _zz__zz__6_14_inner_macOut = ($signed(io_mulInput) * $signed(_6_14_inner_activation));
  assign _zz__zz__6_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_14_inner_macOut)) ? 16'h007f : _zz__6_14_inner_macOut_2);
  assign _zz__6_14_inner_macOut_2 = (($signed(_zz__6_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_14_inner_activation;
    end else begin
      io_macOut = _6_14_inner_macOut;
    end
  end

  assign _zz__6_14_inner_macOut = ($signed(_zz__zz__6_14_inner_macOut) + $signed(_zz__zz__6_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_14_inner_activation <= 8'h00;
      _6_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_14_inner_activation <= io_addInput;
      end else begin
        _6_14_inner_macOut <= _zz__6_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_205 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_13_inner_macOut;
  wire       [15:0]   _zz__zz__6_13_inner_macOut_1;
  wire       [15:0]   _zz__6_13_inner_macOut_1;
  wire       [15:0]   _zz__6_13_inner_macOut_2;
  reg        [7:0]    _6_13_inner_activation;
  reg        [7:0]    _6_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_13_inner_macOut;

  assign _zz__zz__6_13_inner_macOut = ($signed(io_mulInput) * $signed(_6_13_inner_activation));
  assign _zz__zz__6_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_13_inner_macOut)) ? 16'h007f : _zz__6_13_inner_macOut_2);
  assign _zz__6_13_inner_macOut_2 = (($signed(_zz__6_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_13_inner_activation;
    end else begin
      io_macOut = _6_13_inner_macOut;
    end
  end

  assign _zz__6_13_inner_macOut = ($signed(_zz__zz__6_13_inner_macOut) + $signed(_zz__zz__6_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_13_inner_activation <= 8'h00;
      _6_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_13_inner_activation <= io_addInput;
      end else begin
        _6_13_inner_macOut <= _zz__6_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_204 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_12_inner_macOut;
  wire       [15:0]   _zz__zz__6_12_inner_macOut_1;
  wire       [15:0]   _zz__6_12_inner_macOut_1;
  wire       [15:0]   _zz__6_12_inner_macOut_2;
  reg        [7:0]    _6_12_inner_activation;
  reg        [7:0]    _6_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_12_inner_macOut;

  assign _zz__zz__6_12_inner_macOut = ($signed(io_mulInput) * $signed(_6_12_inner_activation));
  assign _zz__zz__6_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_12_inner_macOut)) ? 16'h007f : _zz__6_12_inner_macOut_2);
  assign _zz__6_12_inner_macOut_2 = (($signed(_zz__6_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_12_inner_activation;
    end else begin
      io_macOut = _6_12_inner_macOut;
    end
  end

  assign _zz__6_12_inner_macOut = ($signed(_zz__zz__6_12_inner_macOut) + $signed(_zz__zz__6_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_12_inner_activation <= 8'h00;
      _6_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_12_inner_activation <= io_addInput;
      end else begin
        _6_12_inner_macOut <= _zz__6_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_203 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_11_inner_macOut;
  wire       [15:0]   _zz__zz__6_11_inner_macOut_1;
  wire       [15:0]   _zz__6_11_inner_macOut_1;
  wire       [15:0]   _zz__6_11_inner_macOut_2;
  reg        [7:0]    _6_11_inner_activation;
  reg        [7:0]    _6_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_11_inner_macOut;

  assign _zz__zz__6_11_inner_macOut = ($signed(io_mulInput) * $signed(_6_11_inner_activation));
  assign _zz__zz__6_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_11_inner_macOut)) ? 16'h007f : _zz__6_11_inner_macOut_2);
  assign _zz__6_11_inner_macOut_2 = (($signed(_zz__6_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_11_inner_activation;
    end else begin
      io_macOut = _6_11_inner_macOut;
    end
  end

  assign _zz__6_11_inner_macOut = ($signed(_zz__zz__6_11_inner_macOut) + $signed(_zz__zz__6_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_11_inner_activation <= 8'h00;
      _6_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_11_inner_activation <= io_addInput;
      end else begin
        _6_11_inner_macOut <= _zz__6_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_202 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_10_inner_macOut;
  wire       [15:0]   _zz__zz__6_10_inner_macOut_1;
  wire       [15:0]   _zz__6_10_inner_macOut_1;
  wire       [15:0]   _zz__6_10_inner_macOut_2;
  reg        [7:0]    _6_10_inner_activation;
  reg        [7:0]    _6_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_10_inner_macOut;

  assign _zz__zz__6_10_inner_macOut = ($signed(io_mulInput) * $signed(_6_10_inner_activation));
  assign _zz__zz__6_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_10_inner_macOut)) ? 16'h007f : _zz__6_10_inner_macOut_2);
  assign _zz__6_10_inner_macOut_2 = (($signed(_zz__6_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_10_inner_activation;
    end else begin
      io_macOut = _6_10_inner_macOut;
    end
  end

  assign _zz__6_10_inner_macOut = ($signed(_zz__zz__6_10_inner_macOut) + $signed(_zz__zz__6_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_10_inner_activation <= 8'h00;
      _6_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_10_inner_activation <= io_addInput;
      end else begin
        _6_10_inner_macOut <= _zz__6_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_201 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_9_inner_macOut;
  wire       [15:0]   _zz__zz__6_9_inner_macOut_1;
  wire       [15:0]   _zz__6_9_inner_macOut_1;
  wire       [15:0]   _zz__6_9_inner_macOut_2;
  reg        [7:0]    _6_9_inner_activation;
  reg        [7:0]    _6_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_9_inner_macOut;

  assign _zz__zz__6_9_inner_macOut = ($signed(io_mulInput) * $signed(_6_9_inner_activation));
  assign _zz__zz__6_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_9_inner_macOut)) ? 16'h007f : _zz__6_9_inner_macOut_2);
  assign _zz__6_9_inner_macOut_2 = (($signed(_zz__6_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_9_inner_activation;
    end else begin
      io_macOut = _6_9_inner_macOut;
    end
  end

  assign _zz__6_9_inner_macOut = ($signed(_zz__zz__6_9_inner_macOut) + $signed(_zz__zz__6_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_9_inner_activation <= 8'h00;
      _6_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_9_inner_activation <= io_addInput;
      end else begin
        _6_9_inner_macOut <= _zz__6_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_200 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_8_inner_macOut;
  wire       [15:0]   _zz__zz__6_8_inner_macOut_1;
  wire       [15:0]   _zz__6_8_inner_macOut_1;
  wire       [15:0]   _zz__6_8_inner_macOut_2;
  reg        [7:0]    _6_8_inner_activation;
  reg        [7:0]    _6_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_8_inner_macOut;

  assign _zz__zz__6_8_inner_macOut = ($signed(io_mulInput) * $signed(_6_8_inner_activation));
  assign _zz__zz__6_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_8_inner_macOut)) ? 16'h007f : _zz__6_8_inner_macOut_2);
  assign _zz__6_8_inner_macOut_2 = (($signed(_zz__6_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_8_inner_activation;
    end else begin
      io_macOut = _6_8_inner_macOut;
    end
  end

  assign _zz__6_8_inner_macOut = ($signed(_zz__zz__6_8_inner_macOut) + $signed(_zz__zz__6_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_8_inner_activation <= 8'h00;
      _6_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_8_inner_activation <= io_addInput;
      end else begin
        _6_8_inner_macOut <= _zz__6_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_199 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_7_inner_macOut;
  wire       [15:0]   _zz__zz__6_7_inner_macOut_1;
  wire       [15:0]   _zz__6_7_inner_macOut_1;
  wire       [15:0]   _zz__6_7_inner_macOut_2;
  reg        [7:0]    _6_7_inner_activation;
  reg        [7:0]    _6_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_7_inner_macOut;

  assign _zz__zz__6_7_inner_macOut = ($signed(io_mulInput) * $signed(_6_7_inner_activation));
  assign _zz__zz__6_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_7_inner_macOut)) ? 16'h007f : _zz__6_7_inner_macOut_2);
  assign _zz__6_7_inner_macOut_2 = (($signed(_zz__6_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_7_inner_activation;
    end else begin
      io_macOut = _6_7_inner_macOut;
    end
  end

  assign _zz__6_7_inner_macOut = ($signed(_zz__zz__6_7_inner_macOut) + $signed(_zz__zz__6_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_7_inner_activation <= 8'h00;
      _6_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_7_inner_activation <= io_addInput;
      end else begin
        _6_7_inner_macOut <= _zz__6_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_198 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_6_inner_macOut;
  wire       [15:0]   _zz__zz__6_6_inner_macOut_1;
  wire       [15:0]   _zz__6_6_inner_macOut_1;
  wire       [15:0]   _zz__6_6_inner_macOut_2;
  reg        [7:0]    _6_6_inner_activation;
  reg        [7:0]    _6_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_6_inner_macOut;

  assign _zz__zz__6_6_inner_macOut = ($signed(io_mulInput) * $signed(_6_6_inner_activation));
  assign _zz__zz__6_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_6_inner_macOut)) ? 16'h007f : _zz__6_6_inner_macOut_2);
  assign _zz__6_6_inner_macOut_2 = (($signed(_zz__6_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_6_inner_activation;
    end else begin
      io_macOut = _6_6_inner_macOut;
    end
  end

  assign _zz__6_6_inner_macOut = ($signed(_zz__zz__6_6_inner_macOut) + $signed(_zz__zz__6_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_6_inner_activation <= 8'h00;
      _6_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_6_inner_activation <= io_addInput;
      end else begin
        _6_6_inner_macOut <= _zz__6_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_197 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_5_inner_macOut;
  wire       [15:0]   _zz__zz__6_5_inner_macOut_1;
  wire       [15:0]   _zz__6_5_inner_macOut_1;
  wire       [15:0]   _zz__6_5_inner_macOut_2;
  reg        [7:0]    _6_5_inner_activation;
  reg        [7:0]    _6_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_5_inner_macOut;

  assign _zz__zz__6_5_inner_macOut = ($signed(io_mulInput) * $signed(_6_5_inner_activation));
  assign _zz__zz__6_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_5_inner_macOut)) ? 16'h007f : _zz__6_5_inner_macOut_2);
  assign _zz__6_5_inner_macOut_2 = (($signed(_zz__6_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_5_inner_activation;
    end else begin
      io_macOut = _6_5_inner_macOut;
    end
  end

  assign _zz__6_5_inner_macOut = ($signed(_zz__zz__6_5_inner_macOut) + $signed(_zz__zz__6_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_5_inner_activation <= 8'h00;
      _6_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_5_inner_activation <= io_addInput;
      end else begin
        _6_5_inner_macOut <= _zz__6_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_196 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_4_inner_macOut;
  wire       [15:0]   _zz__zz__6_4_inner_macOut_1;
  wire       [15:0]   _zz__6_4_inner_macOut_1;
  wire       [15:0]   _zz__6_4_inner_macOut_2;
  reg        [7:0]    _6_4_inner_activation;
  reg        [7:0]    _6_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_4_inner_macOut;

  assign _zz__zz__6_4_inner_macOut = ($signed(io_mulInput) * $signed(_6_4_inner_activation));
  assign _zz__zz__6_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_4_inner_macOut)) ? 16'h007f : _zz__6_4_inner_macOut_2);
  assign _zz__6_4_inner_macOut_2 = (($signed(_zz__6_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_4_inner_activation;
    end else begin
      io_macOut = _6_4_inner_macOut;
    end
  end

  assign _zz__6_4_inner_macOut = ($signed(_zz__zz__6_4_inner_macOut) + $signed(_zz__zz__6_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_4_inner_activation <= 8'h00;
      _6_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_4_inner_activation <= io_addInput;
      end else begin
        _6_4_inner_macOut <= _zz__6_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_195 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_3_inner_macOut;
  wire       [15:0]   _zz__zz__6_3_inner_macOut_1;
  wire       [15:0]   _zz__6_3_inner_macOut_1;
  wire       [15:0]   _zz__6_3_inner_macOut_2;
  reg        [7:0]    _6_3_inner_activation;
  reg        [7:0]    _6_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_3_inner_macOut;

  assign _zz__zz__6_3_inner_macOut = ($signed(io_mulInput) * $signed(_6_3_inner_activation));
  assign _zz__zz__6_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_3_inner_macOut)) ? 16'h007f : _zz__6_3_inner_macOut_2);
  assign _zz__6_3_inner_macOut_2 = (($signed(_zz__6_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_3_inner_activation;
    end else begin
      io_macOut = _6_3_inner_macOut;
    end
  end

  assign _zz__6_3_inner_macOut = ($signed(_zz__zz__6_3_inner_macOut) + $signed(_zz__zz__6_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_3_inner_activation <= 8'h00;
      _6_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_3_inner_activation <= io_addInput;
      end else begin
        _6_3_inner_macOut <= _zz__6_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_194 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_2_inner_macOut;
  wire       [15:0]   _zz__zz__6_2_inner_macOut_1;
  wire       [15:0]   _zz__6_2_inner_macOut_1;
  wire       [15:0]   _zz__6_2_inner_macOut_2;
  reg        [7:0]    _6_2_inner_activation;
  reg        [7:0]    _6_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_2_inner_macOut;

  assign _zz__zz__6_2_inner_macOut = ($signed(io_mulInput) * $signed(_6_2_inner_activation));
  assign _zz__zz__6_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_2_inner_macOut)) ? 16'h007f : _zz__6_2_inner_macOut_2);
  assign _zz__6_2_inner_macOut_2 = (($signed(_zz__6_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_2_inner_activation;
    end else begin
      io_macOut = _6_2_inner_macOut;
    end
  end

  assign _zz__6_2_inner_macOut = ($signed(_zz__zz__6_2_inner_macOut) + $signed(_zz__zz__6_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_2_inner_activation <= 8'h00;
      _6_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_2_inner_activation <= io_addInput;
      end else begin
        _6_2_inner_macOut <= _zz__6_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_193 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_1_inner_macOut;
  wire       [15:0]   _zz__zz__6_1_inner_macOut_1;
  wire       [15:0]   _zz__6_1_inner_macOut_1;
  wire       [15:0]   _zz__6_1_inner_macOut_2;
  reg        [7:0]    _6_1_inner_activation;
  reg        [7:0]    _6_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_1_inner_macOut;

  assign _zz__zz__6_1_inner_macOut = ($signed(io_mulInput) * $signed(_6_1_inner_activation));
  assign _zz__zz__6_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_1_inner_macOut)) ? 16'h007f : _zz__6_1_inner_macOut_2);
  assign _zz__6_1_inner_macOut_2 = (($signed(_zz__6_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_1_inner_activation;
    end else begin
      io_macOut = _6_1_inner_macOut;
    end
  end

  assign _zz__6_1_inner_macOut = ($signed(_zz__zz__6_1_inner_macOut) + $signed(_zz__zz__6_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_1_inner_activation <= 8'h00;
      _6_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_1_inner_activation <= io_addInput;
      end else begin
        _6_1_inner_macOut <= _zz__6_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_192 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__6_0_inner_macOut;
  wire       [15:0]   _zz__zz__6_0_inner_macOut_1;
  wire       [15:0]   _zz__6_0_inner_macOut_1;
  wire       [15:0]   _zz__6_0_inner_macOut_2;
  reg        [7:0]    _6_0_inner_activation;
  reg        [7:0]    _6_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__6_0_inner_macOut;

  assign _zz__zz__6_0_inner_macOut = ($signed(io_mulInput) * $signed(_6_0_inner_activation));
  assign _zz__zz__6_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__6_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__6_0_inner_macOut)) ? 16'h007f : _zz__6_0_inner_macOut_2);
  assign _zz__6_0_inner_macOut_2 = (($signed(_zz__6_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__6_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _6_0_inner_activation;
    end else begin
      io_macOut = _6_0_inner_macOut;
    end
  end

  assign _zz__6_0_inner_macOut = ($signed(_zz__zz__6_0_inner_macOut) + $signed(_zz__zz__6_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _6_0_inner_activation <= 8'h00;
      _6_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _6_0_inner_activation <= io_addInput;
      end else begin
        _6_0_inner_macOut <= _zz__6_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_191 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_31_inner_macOut;
  wire       [15:0]   _zz__zz__5_31_inner_macOut_1;
  wire       [15:0]   _zz__5_31_inner_macOut_1;
  wire       [15:0]   _zz__5_31_inner_macOut_2;
  reg        [7:0]    _5_31_inner_activation;
  reg        [7:0]    _5_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_31_inner_macOut;

  assign _zz__zz__5_31_inner_macOut = ($signed(io_mulInput) * $signed(_5_31_inner_activation));
  assign _zz__zz__5_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_31_inner_macOut)) ? 16'h007f : _zz__5_31_inner_macOut_2);
  assign _zz__5_31_inner_macOut_2 = (($signed(_zz__5_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_31_inner_activation;
    end else begin
      io_macOut = _5_31_inner_macOut;
    end
  end

  assign _zz__5_31_inner_macOut = ($signed(_zz__zz__5_31_inner_macOut) + $signed(_zz__zz__5_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_31_inner_activation <= 8'h00;
      _5_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_31_inner_activation <= io_addInput;
      end else begin
        _5_31_inner_macOut <= _zz__5_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_190 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_30_inner_macOut;
  wire       [15:0]   _zz__zz__5_30_inner_macOut_1;
  wire       [15:0]   _zz__5_30_inner_macOut_1;
  wire       [15:0]   _zz__5_30_inner_macOut_2;
  reg        [7:0]    _5_30_inner_activation;
  reg        [7:0]    _5_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_30_inner_macOut;

  assign _zz__zz__5_30_inner_macOut = ($signed(io_mulInput) * $signed(_5_30_inner_activation));
  assign _zz__zz__5_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_30_inner_macOut)) ? 16'h007f : _zz__5_30_inner_macOut_2);
  assign _zz__5_30_inner_macOut_2 = (($signed(_zz__5_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_30_inner_activation;
    end else begin
      io_macOut = _5_30_inner_macOut;
    end
  end

  assign _zz__5_30_inner_macOut = ($signed(_zz__zz__5_30_inner_macOut) + $signed(_zz__zz__5_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_30_inner_activation <= 8'h00;
      _5_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_30_inner_activation <= io_addInput;
      end else begin
        _5_30_inner_macOut <= _zz__5_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_189 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_29_inner_macOut;
  wire       [15:0]   _zz__zz__5_29_inner_macOut_1;
  wire       [15:0]   _zz__5_29_inner_macOut_1;
  wire       [15:0]   _zz__5_29_inner_macOut_2;
  reg        [7:0]    _5_29_inner_activation;
  reg        [7:0]    _5_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_29_inner_macOut;

  assign _zz__zz__5_29_inner_macOut = ($signed(io_mulInput) * $signed(_5_29_inner_activation));
  assign _zz__zz__5_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_29_inner_macOut)) ? 16'h007f : _zz__5_29_inner_macOut_2);
  assign _zz__5_29_inner_macOut_2 = (($signed(_zz__5_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_29_inner_activation;
    end else begin
      io_macOut = _5_29_inner_macOut;
    end
  end

  assign _zz__5_29_inner_macOut = ($signed(_zz__zz__5_29_inner_macOut) + $signed(_zz__zz__5_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_29_inner_activation <= 8'h00;
      _5_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_29_inner_activation <= io_addInput;
      end else begin
        _5_29_inner_macOut <= _zz__5_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_188 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_28_inner_macOut;
  wire       [15:0]   _zz__zz__5_28_inner_macOut_1;
  wire       [15:0]   _zz__5_28_inner_macOut_1;
  wire       [15:0]   _zz__5_28_inner_macOut_2;
  reg        [7:0]    _5_28_inner_activation;
  reg        [7:0]    _5_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_28_inner_macOut;

  assign _zz__zz__5_28_inner_macOut = ($signed(io_mulInput) * $signed(_5_28_inner_activation));
  assign _zz__zz__5_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_28_inner_macOut)) ? 16'h007f : _zz__5_28_inner_macOut_2);
  assign _zz__5_28_inner_macOut_2 = (($signed(_zz__5_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_28_inner_activation;
    end else begin
      io_macOut = _5_28_inner_macOut;
    end
  end

  assign _zz__5_28_inner_macOut = ($signed(_zz__zz__5_28_inner_macOut) + $signed(_zz__zz__5_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_28_inner_activation <= 8'h00;
      _5_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_28_inner_activation <= io_addInput;
      end else begin
        _5_28_inner_macOut <= _zz__5_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_187 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_27_inner_macOut;
  wire       [15:0]   _zz__zz__5_27_inner_macOut_1;
  wire       [15:0]   _zz__5_27_inner_macOut_1;
  wire       [15:0]   _zz__5_27_inner_macOut_2;
  reg        [7:0]    _5_27_inner_activation;
  reg        [7:0]    _5_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_27_inner_macOut;

  assign _zz__zz__5_27_inner_macOut = ($signed(io_mulInput) * $signed(_5_27_inner_activation));
  assign _zz__zz__5_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_27_inner_macOut)) ? 16'h007f : _zz__5_27_inner_macOut_2);
  assign _zz__5_27_inner_macOut_2 = (($signed(_zz__5_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_27_inner_activation;
    end else begin
      io_macOut = _5_27_inner_macOut;
    end
  end

  assign _zz__5_27_inner_macOut = ($signed(_zz__zz__5_27_inner_macOut) + $signed(_zz__zz__5_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_27_inner_activation <= 8'h00;
      _5_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_27_inner_activation <= io_addInput;
      end else begin
        _5_27_inner_macOut <= _zz__5_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_186 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_26_inner_macOut;
  wire       [15:0]   _zz__zz__5_26_inner_macOut_1;
  wire       [15:0]   _zz__5_26_inner_macOut_1;
  wire       [15:0]   _zz__5_26_inner_macOut_2;
  reg        [7:0]    _5_26_inner_activation;
  reg        [7:0]    _5_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_26_inner_macOut;

  assign _zz__zz__5_26_inner_macOut = ($signed(io_mulInput) * $signed(_5_26_inner_activation));
  assign _zz__zz__5_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_26_inner_macOut)) ? 16'h007f : _zz__5_26_inner_macOut_2);
  assign _zz__5_26_inner_macOut_2 = (($signed(_zz__5_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_26_inner_activation;
    end else begin
      io_macOut = _5_26_inner_macOut;
    end
  end

  assign _zz__5_26_inner_macOut = ($signed(_zz__zz__5_26_inner_macOut) + $signed(_zz__zz__5_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_26_inner_activation <= 8'h00;
      _5_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_26_inner_activation <= io_addInput;
      end else begin
        _5_26_inner_macOut <= _zz__5_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_185 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_25_inner_macOut;
  wire       [15:0]   _zz__zz__5_25_inner_macOut_1;
  wire       [15:0]   _zz__5_25_inner_macOut_1;
  wire       [15:0]   _zz__5_25_inner_macOut_2;
  reg        [7:0]    _5_25_inner_activation;
  reg        [7:0]    _5_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_25_inner_macOut;

  assign _zz__zz__5_25_inner_macOut = ($signed(io_mulInput) * $signed(_5_25_inner_activation));
  assign _zz__zz__5_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_25_inner_macOut)) ? 16'h007f : _zz__5_25_inner_macOut_2);
  assign _zz__5_25_inner_macOut_2 = (($signed(_zz__5_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_25_inner_activation;
    end else begin
      io_macOut = _5_25_inner_macOut;
    end
  end

  assign _zz__5_25_inner_macOut = ($signed(_zz__zz__5_25_inner_macOut) + $signed(_zz__zz__5_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_25_inner_activation <= 8'h00;
      _5_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_25_inner_activation <= io_addInput;
      end else begin
        _5_25_inner_macOut <= _zz__5_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_184 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_24_inner_macOut;
  wire       [15:0]   _zz__zz__5_24_inner_macOut_1;
  wire       [15:0]   _zz__5_24_inner_macOut_1;
  wire       [15:0]   _zz__5_24_inner_macOut_2;
  reg        [7:0]    _5_24_inner_activation;
  reg        [7:0]    _5_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_24_inner_macOut;

  assign _zz__zz__5_24_inner_macOut = ($signed(io_mulInput) * $signed(_5_24_inner_activation));
  assign _zz__zz__5_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_24_inner_macOut)) ? 16'h007f : _zz__5_24_inner_macOut_2);
  assign _zz__5_24_inner_macOut_2 = (($signed(_zz__5_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_24_inner_activation;
    end else begin
      io_macOut = _5_24_inner_macOut;
    end
  end

  assign _zz__5_24_inner_macOut = ($signed(_zz__zz__5_24_inner_macOut) + $signed(_zz__zz__5_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_24_inner_activation <= 8'h00;
      _5_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_24_inner_activation <= io_addInput;
      end else begin
        _5_24_inner_macOut <= _zz__5_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_183 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_23_inner_macOut;
  wire       [15:0]   _zz__zz__5_23_inner_macOut_1;
  wire       [15:0]   _zz__5_23_inner_macOut_1;
  wire       [15:0]   _zz__5_23_inner_macOut_2;
  reg        [7:0]    _5_23_inner_activation;
  reg        [7:0]    _5_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_23_inner_macOut;

  assign _zz__zz__5_23_inner_macOut = ($signed(io_mulInput) * $signed(_5_23_inner_activation));
  assign _zz__zz__5_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_23_inner_macOut)) ? 16'h007f : _zz__5_23_inner_macOut_2);
  assign _zz__5_23_inner_macOut_2 = (($signed(_zz__5_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_23_inner_activation;
    end else begin
      io_macOut = _5_23_inner_macOut;
    end
  end

  assign _zz__5_23_inner_macOut = ($signed(_zz__zz__5_23_inner_macOut) + $signed(_zz__zz__5_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_23_inner_activation <= 8'h00;
      _5_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_23_inner_activation <= io_addInput;
      end else begin
        _5_23_inner_macOut <= _zz__5_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_182 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_22_inner_macOut;
  wire       [15:0]   _zz__zz__5_22_inner_macOut_1;
  wire       [15:0]   _zz__5_22_inner_macOut_1;
  wire       [15:0]   _zz__5_22_inner_macOut_2;
  reg        [7:0]    _5_22_inner_activation;
  reg        [7:0]    _5_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_22_inner_macOut;

  assign _zz__zz__5_22_inner_macOut = ($signed(io_mulInput) * $signed(_5_22_inner_activation));
  assign _zz__zz__5_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_22_inner_macOut)) ? 16'h007f : _zz__5_22_inner_macOut_2);
  assign _zz__5_22_inner_macOut_2 = (($signed(_zz__5_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_22_inner_activation;
    end else begin
      io_macOut = _5_22_inner_macOut;
    end
  end

  assign _zz__5_22_inner_macOut = ($signed(_zz__zz__5_22_inner_macOut) + $signed(_zz__zz__5_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_22_inner_activation <= 8'h00;
      _5_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_22_inner_activation <= io_addInput;
      end else begin
        _5_22_inner_macOut <= _zz__5_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_181 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_21_inner_macOut;
  wire       [15:0]   _zz__zz__5_21_inner_macOut_1;
  wire       [15:0]   _zz__5_21_inner_macOut_1;
  wire       [15:0]   _zz__5_21_inner_macOut_2;
  reg        [7:0]    _5_21_inner_activation;
  reg        [7:0]    _5_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_21_inner_macOut;

  assign _zz__zz__5_21_inner_macOut = ($signed(io_mulInput) * $signed(_5_21_inner_activation));
  assign _zz__zz__5_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_21_inner_macOut)) ? 16'h007f : _zz__5_21_inner_macOut_2);
  assign _zz__5_21_inner_macOut_2 = (($signed(_zz__5_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_21_inner_activation;
    end else begin
      io_macOut = _5_21_inner_macOut;
    end
  end

  assign _zz__5_21_inner_macOut = ($signed(_zz__zz__5_21_inner_macOut) + $signed(_zz__zz__5_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_21_inner_activation <= 8'h00;
      _5_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_21_inner_activation <= io_addInput;
      end else begin
        _5_21_inner_macOut <= _zz__5_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_180 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_20_inner_macOut;
  wire       [15:0]   _zz__zz__5_20_inner_macOut_1;
  wire       [15:0]   _zz__5_20_inner_macOut_1;
  wire       [15:0]   _zz__5_20_inner_macOut_2;
  reg        [7:0]    _5_20_inner_activation;
  reg        [7:0]    _5_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_20_inner_macOut;

  assign _zz__zz__5_20_inner_macOut = ($signed(io_mulInput) * $signed(_5_20_inner_activation));
  assign _zz__zz__5_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_20_inner_macOut)) ? 16'h007f : _zz__5_20_inner_macOut_2);
  assign _zz__5_20_inner_macOut_2 = (($signed(_zz__5_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_20_inner_activation;
    end else begin
      io_macOut = _5_20_inner_macOut;
    end
  end

  assign _zz__5_20_inner_macOut = ($signed(_zz__zz__5_20_inner_macOut) + $signed(_zz__zz__5_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_20_inner_activation <= 8'h00;
      _5_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_20_inner_activation <= io_addInput;
      end else begin
        _5_20_inner_macOut <= _zz__5_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_179 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_19_inner_macOut;
  wire       [15:0]   _zz__zz__5_19_inner_macOut_1;
  wire       [15:0]   _zz__5_19_inner_macOut_1;
  wire       [15:0]   _zz__5_19_inner_macOut_2;
  reg        [7:0]    _5_19_inner_activation;
  reg        [7:0]    _5_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_19_inner_macOut;

  assign _zz__zz__5_19_inner_macOut = ($signed(io_mulInput) * $signed(_5_19_inner_activation));
  assign _zz__zz__5_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_19_inner_macOut)) ? 16'h007f : _zz__5_19_inner_macOut_2);
  assign _zz__5_19_inner_macOut_2 = (($signed(_zz__5_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_19_inner_activation;
    end else begin
      io_macOut = _5_19_inner_macOut;
    end
  end

  assign _zz__5_19_inner_macOut = ($signed(_zz__zz__5_19_inner_macOut) + $signed(_zz__zz__5_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_19_inner_activation <= 8'h00;
      _5_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_19_inner_activation <= io_addInput;
      end else begin
        _5_19_inner_macOut <= _zz__5_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_178 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_18_inner_macOut;
  wire       [15:0]   _zz__zz__5_18_inner_macOut_1;
  wire       [15:0]   _zz__5_18_inner_macOut_1;
  wire       [15:0]   _zz__5_18_inner_macOut_2;
  reg        [7:0]    _5_18_inner_activation;
  reg        [7:0]    _5_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_18_inner_macOut;

  assign _zz__zz__5_18_inner_macOut = ($signed(io_mulInput) * $signed(_5_18_inner_activation));
  assign _zz__zz__5_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_18_inner_macOut)) ? 16'h007f : _zz__5_18_inner_macOut_2);
  assign _zz__5_18_inner_macOut_2 = (($signed(_zz__5_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_18_inner_activation;
    end else begin
      io_macOut = _5_18_inner_macOut;
    end
  end

  assign _zz__5_18_inner_macOut = ($signed(_zz__zz__5_18_inner_macOut) + $signed(_zz__zz__5_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_18_inner_activation <= 8'h00;
      _5_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_18_inner_activation <= io_addInput;
      end else begin
        _5_18_inner_macOut <= _zz__5_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_177 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_17_inner_macOut;
  wire       [15:0]   _zz__zz__5_17_inner_macOut_1;
  wire       [15:0]   _zz__5_17_inner_macOut_1;
  wire       [15:0]   _zz__5_17_inner_macOut_2;
  reg        [7:0]    _5_17_inner_activation;
  reg        [7:0]    _5_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_17_inner_macOut;

  assign _zz__zz__5_17_inner_macOut = ($signed(io_mulInput) * $signed(_5_17_inner_activation));
  assign _zz__zz__5_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_17_inner_macOut)) ? 16'h007f : _zz__5_17_inner_macOut_2);
  assign _zz__5_17_inner_macOut_2 = (($signed(_zz__5_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_17_inner_activation;
    end else begin
      io_macOut = _5_17_inner_macOut;
    end
  end

  assign _zz__5_17_inner_macOut = ($signed(_zz__zz__5_17_inner_macOut) + $signed(_zz__zz__5_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_17_inner_activation <= 8'h00;
      _5_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_17_inner_activation <= io_addInput;
      end else begin
        _5_17_inner_macOut <= _zz__5_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_176 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_16_inner_macOut;
  wire       [15:0]   _zz__zz__5_16_inner_macOut_1;
  wire       [15:0]   _zz__5_16_inner_macOut_1;
  wire       [15:0]   _zz__5_16_inner_macOut_2;
  reg        [7:0]    _5_16_inner_activation;
  reg        [7:0]    _5_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_16_inner_macOut;

  assign _zz__zz__5_16_inner_macOut = ($signed(io_mulInput) * $signed(_5_16_inner_activation));
  assign _zz__zz__5_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_16_inner_macOut)) ? 16'h007f : _zz__5_16_inner_macOut_2);
  assign _zz__5_16_inner_macOut_2 = (($signed(_zz__5_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_16_inner_activation;
    end else begin
      io_macOut = _5_16_inner_macOut;
    end
  end

  assign _zz__5_16_inner_macOut = ($signed(_zz__zz__5_16_inner_macOut) + $signed(_zz__zz__5_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_16_inner_activation <= 8'h00;
      _5_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_16_inner_activation <= io_addInput;
      end else begin
        _5_16_inner_macOut <= _zz__5_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_175 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_15_inner_macOut;
  wire       [15:0]   _zz__zz__5_15_inner_macOut_1;
  wire       [15:0]   _zz__5_15_inner_macOut_1;
  wire       [15:0]   _zz__5_15_inner_macOut_2;
  reg        [7:0]    _5_15_inner_activation;
  reg        [7:0]    _5_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_15_inner_macOut;

  assign _zz__zz__5_15_inner_macOut = ($signed(io_mulInput) * $signed(_5_15_inner_activation));
  assign _zz__zz__5_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_15_inner_macOut)) ? 16'h007f : _zz__5_15_inner_macOut_2);
  assign _zz__5_15_inner_macOut_2 = (($signed(_zz__5_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_15_inner_activation;
    end else begin
      io_macOut = _5_15_inner_macOut;
    end
  end

  assign _zz__5_15_inner_macOut = ($signed(_zz__zz__5_15_inner_macOut) + $signed(_zz__zz__5_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_15_inner_activation <= 8'h00;
      _5_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_15_inner_activation <= io_addInput;
      end else begin
        _5_15_inner_macOut <= _zz__5_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_174 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_14_inner_macOut;
  wire       [15:0]   _zz__zz__5_14_inner_macOut_1;
  wire       [15:0]   _zz__5_14_inner_macOut_1;
  wire       [15:0]   _zz__5_14_inner_macOut_2;
  reg        [7:0]    _5_14_inner_activation;
  reg        [7:0]    _5_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_14_inner_macOut;

  assign _zz__zz__5_14_inner_macOut = ($signed(io_mulInput) * $signed(_5_14_inner_activation));
  assign _zz__zz__5_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_14_inner_macOut)) ? 16'h007f : _zz__5_14_inner_macOut_2);
  assign _zz__5_14_inner_macOut_2 = (($signed(_zz__5_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_14_inner_activation;
    end else begin
      io_macOut = _5_14_inner_macOut;
    end
  end

  assign _zz__5_14_inner_macOut = ($signed(_zz__zz__5_14_inner_macOut) + $signed(_zz__zz__5_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_14_inner_activation <= 8'h00;
      _5_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_14_inner_activation <= io_addInput;
      end else begin
        _5_14_inner_macOut <= _zz__5_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_173 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_13_inner_macOut;
  wire       [15:0]   _zz__zz__5_13_inner_macOut_1;
  wire       [15:0]   _zz__5_13_inner_macOut_1;
  wire       [15:0]   _zz__5_13_inner_macOut_2;
  reg        [7:0]    _5_13_inner_activation;
  reg        [7:0]    _5_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_13_inner_macOut;

  assign _zz__zz__5_13_inner_macOut = ($signed(io_mulInput) * $signed(_5_13_inner_activation));
  assign _zz__zz__5_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_13_inner_macOut)) ? 16'h007f : _zz__5_13_inner_macOut_2);
  assign _zz__5_13_inner_macOut_2 = (($signed(_zz__5_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_13_inner_activation;
    end else begin
      io_macOut = _5_13_inner_macOut;
    end
  end

  assign _zz__5_13_inner_macOut = ($signed(_zz__zz__5_13_inner_macOut) + $signed(_zz__zz__5_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_13_inner_activation <= 8'h00;
      _5_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_13_inner_activation <= io_addInput;
      end else begin
        _5_13_inner_macOut <= _zz__5_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_172 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_12_inner_macOut;
  wire       [15:0]   _zz__zz__5_12_inner_macOut_1;
  wire       [15:0]   _zz__5_12_inner_macOut_1;
  wire       [15:0]   _zz__5_12_inner_macOut_2;
  reg        [7:0]    _5_12_inner_activation;
  reg        [7:0]    _5_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_12_inner_macOut;

  assign _zz__zz__5_12_inner_macOut = ($signed(io_mulInput) * $signed(_5_12_inner_activation));
  assign _zz__zz__5_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_12_inner_macOut)) ? 16'h007f : _zz__5_12_inner_macOut_2);
  assign _zz__5_12_inner_macOut_2 = (($signed(_zz__5_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_12_inner_activation;
    end else begin
      io_macOut = _5_12_inner_macOut;
    end
  end

  assign _zz__5_12_inner_macOut = ($signed(_zz__zz__5_12_inner_macOut) + $signed(_zz__zz__5_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_12_inner_activation <= 8'h00;
      _5_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_12_inner_activation <= io_addInput;
      end else begin
        _5_12_inner_macOut <= _zz__5_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_171 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_11_inner_macOut;
  wire       [15:0]   _zz__zz__5_11_inner_macOut_1;
  wire       [15:0]   _zz__5_11_inner_macOut_1;
  wire       [15:0]   _zz__5_11_inner_macOut_2;
  reg        [7:0]    _5_11_inner_activation;
  reg        [7:0]    _5_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_11_inner_macOut;

  assign _zz__zz__5_11_inner_macOut = ($signed(io_mulInput) * $signed(_5_11_inner_activation));
  assign _zz__zz__5_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_11_inner_macOut)) ? 16'h007f : _zz__5_11_inner_macOut_2);
  assign _zz__5_11_inner_macOut_2 = (($signed(_zz__5_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_11_inner_activation;
    end else begin
      io_macOut = _5_11_inner_macOut;
    end
  end

  assign _zz__5_11_inner_macOut = ($signed(_zz__zz__5_11_inner_macOut) + $signed(_zz__zz__5_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_11_inner_activation <= 8'h00;
      _5_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_11_inner_activation <= io_addInput;
      end else begin
        _5_11_inner_macOut <= _zz__5_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_170 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_10_inner_macOut;
  wire       [15:0]   _zz__zz__5_10_inner_macOut_1;
  wire       [15:0]   _zz__5_10_inner_macOut_1;
  wire       [15:0]   _zz__5_10_inner_macOut_2;
  reg        [7:0]    _5_10_inner_activation;
  reg        [7:0]    _5_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_10_inner_macOut;

  assign _zz__zz__5_10_inner_macOut = ($signed(io_mulInput) * $signed(_5_10_inner_activation));
  assign _zz__zz__5_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_10_inner_macOut)) ? 16'h007f : _zz__5_10_inner_macOut_2);
  assign _zz__5_10_inner_macOut_2 = (($signed(_zz__5_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_10_inner_activation;
    end else begin
      io_macOut = _5_10_inner_macOut;
    end
  end

  assign _zz__5_10_inner_macOut = ($signed(_zz__zz__5_10_inner_macOut) + $signed(_zz__zz__5_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_10_inner_activation <= 8'h00;
      _5_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_10_inner_activation <= io_addInput;
      end else begin
        _5_10_inner_macOut <= _zz__5_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_169 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_9_inner_macOut;
  wire       [15:0]   _zz__zz__5_9_inner_macOut_1;
  wire       [15:0]   _zz__5_9_inner_macOut_1;
  wire       [15:0]   _zz__5_9_inner_macOut_2;
  reg        [7:0]    _5_9_inner_activation;
  reg        [7:0]    _5_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_9_inner_macOut;

  assign _zz__zz__5_9_inner_macOut = ($signed(io_mulInput) * $signed(_5_9_inner_activation));
  assign _zz__zz__5_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_9_inner_macOut)) ? 16'h007f : _zz__5_9_inner_macOut_2);
  assign _zz__5_9_inner_macOut_2 = (($signed(_zz__5_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_9_inner_activation;
    end else begin
      io_macOut = _5_9_inner_macOut;
    end
  end

  assign _zz__5_9_inner_macOut = ($signed(_zz__zz__5_9_inner_macOut) + $signed(_zz__zz__5_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_9_inner_activation <= 8'h00;
      _5_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_9_inner_activation <= io_addInput;
      end else begin
        _5_9_inner_macOut <= _zz__5_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_168 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_8_inner_macOut;
  wire       [15:0]   _zz__zz__5_8_inner_macOut_1;
  wire       [15:0]   _zz__5_8_inner_macOut_1;
  wire       [15:0]   _zz__5_8_inner_macOut_2;
  reg        [7:0]    _5_8_inner_activation;
  reg        [7:0]    _5_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_8_inner_macOut;

  assign _zz__zz__5_8_inner_macOut = ($signed(io_mulInput) * $signed(_5_8_inner_activation));
  assign _zz__zz__5_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_8_inner_macOut)) ? 16'h007f : _zz__5_8_inner_macOut_2);
  assign _zz__5_8_inner_macOut_2 = (($signed(_zz__5_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_8_inner_activation;
    end else begin
      io_macOut = _5_8_inner_macOut;
    end
  end

  assign _zz__5_8_inner_macOut = ($signed(_zz__zz__5_8_inner_macOut) + $signed(_zz__zz__5_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_8_inner_activation <= 8'h00;
      _5_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_8_inner_activation <= io_addInput;
      end else begin
        _5_8_inner_macOut <= _zz__5_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_167 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_7_inner_macOut;
  wire       [15:0]   _zz__zz__5_7_inner_macOut_1;
  wire       [15:0]   _zz__5_7_inner_macOut_1;
  wire       [15:0]   _zz__5_7_inner_macOut_2;
  reg        [7:0]    _5_7_inner_activation;
  reg        [7:0]    _5_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_7_inner_macOut;

  assign _zz__zz__5_7_inner_macOut = ($signed(io_mulInput) * $signed(_5_7_inner_activation));
  assign _zz__zz__5_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_7_inner_macOut)) ? 16'h007f : _zz__5_7_inner_macOut_2);
  assign _zz__5_7_inner_macOut_2 = (($signed(_zz__5_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_7_inner_activation;
    end else begin
      io_macOut = _5_7_inner_macOut;
    end
  end

  assign _zz__5_7_inner_macOut = ($signed(_zz__zz__5_7_inner_macOut) + $signed(_zz__zz__5_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_7_inner_activation <= 8'h00;
      _5_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_7_inner_activation <= io_addInput;
      end else begin
        _5_7_inner_macOut <= _zz__5_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_166 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_6_inner_macOut;
  wire       [15:0]   _zz__zz__5_6_inner_macOut_1;
  wire       [15:0]   _zz__5_6_inner_macOut_1;
  wire       [15:0]   _zz__5_6_inner_macOut_2;
  reg        [7:0]    _5_6_inner_activation;
  reg        [7:0]    _5_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_6_inner_macOut;

  assign _zz__zz__5_6_inner_macOut = ($signed(io_mulInput) * $signed(_5_6_inner_activation));
  assign _zz__zz__5_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_6_inner_macOut)) ? 16'h007f : _zz__5_6_inner_macOut_2);
  assign _zz__5_6_inner_macOut_2 = (($signed(_zz__5_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_6_inner_activation;
    end else begin
      io_macOut = _5_6_inner_macOut;
    end
  end

  assign _zz__5_6_inner_macOut = ($signed(_zz__zz__5_6_inner_macOut) + $signed(_zz__zz__5_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_6_inner_activation <= 8'h00;
      _5_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_6_inner_activation <= io_addInput;
      end else begin
        _5_6_inner_macOut <= _zz__5_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_165 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_5_inner_macOut;
  wire       [15:0]   _zz__zz__5_5_inner_macOut_1;
  wire       [15:0]   _zz__5_5_inner_macOut_1;
  wire       [15:0]   _zz__5_5_inner_macOut_2;
  reg        [7:0]    _5_5_inner_activation;
  reg        [7:0]    _5_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_5_inner_macOut;

  assign _zz__zz__5_5_inner_macOut = ($signed(io_mulInput) * $signed(_5_5_inner_activation));
  assign _zz__zz__5_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_5_inner_macOut)) ? 16'h007f : _zz__5_5_inner_macOut_2);
  assign _zz__5_5_inner_macOut_2 = (($signed(_zz__5_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_5_inner_activation;
    end else begin
      io_macOut = _5_5_inner_macOut;
    end
  end

  assign _zz__5_5_inner_macOut = ($signed(_zz__zz__5_5_inner_macOut) + $signed(_zz__zz__5_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_5_inner_activation <= 8'h00;
      _5_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_5_inner_activation <= io_addInput;
      end else begin
        _5_5_inner_macOut <= _zz__5_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_164 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_4_inner_macOut;
  wire       [15:0]   _zz__zz__5_4_inner_macOut_1;
  wire       [15:0]   _zz__5_4_inner_macOut_1;
  wire       [15:0]   _zz__5_4_inner_macOut_2;
  reg        [7:0]    _5_4_inner_activation;
  reg        [7:0]    _5_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_4_inner_macOut;

  assign _zz__zz__5_4_inner_macOut = ($signed(io_mulInput) * $signed(_5_4_inner_activation));
  assign _zz__zz__5_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_4_inner_macOut)) ? 16'h007f : _zz__5_4_inner_macOut_2);
  assign _zz__5_4_inner_macOut_2 = (($signed(_zz__5_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_4_inner_activation;
    end else begin
      io_macOut = _5_4_inner_macOut;
    end
  end

  assign _zz__5_4_inner_macOut = ($signed(_zz__zz__5_4_inner_macOut) + $signed(_zz__zz__5_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_4_inner_activation <= 8'h00;
      _5_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_4_inner_activation <= io_addInput;
      end else begin
        _5_4_inner_macOut <= _zz__5_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_163 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_3_inner_macOut;
  wire       [15:0]   _zz__zz__5_3_inner_macOut_1;
  wire       [15:0]   _zz__5_3_inner_macOut_1;
  wire       [15:0]   _zz__5_3_inner_macOut_2;
  reg        [7:0]    _5_3_inner_activation;
  reg        [7:0]    _5_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_3_inner_macOut;

  assign _zz__zz__5_3_inner_macOut = ($signed(io_mulInput) * $signed(_5_3_inner_activation));
  assign _zz__zz__5_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_3_inner_macOut)) ? 16'h007f : _zz__5_3_inner_macOut_2);
  assign _zz__5_3_inner_macOut_2 = (($signed(_zz__5_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_3_inner_activation;
    end else begin
      io_macOut = _5_3_inner_macOut;
    end
  end

  assign _zz__5_3_inner_macOut = ($signed(_zz__zz__5_3_inner_macOut) + $signed(_zz__zz__5_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_3_inner_activation <= 8'h00;
      _5_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_3_inner_activation <= io_addInput;
      end else begin
        _5_3_inner_macOut <= _zz__5_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_162 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_2_inner_macOut;
  wire       [15:0]   _zz__zz__5_2_inner_macOut_1;
  wire       [15:0]   _zz__5_2_inner_macOut_1;
  wire       [15:0]   _zz__5_2_inner_macOut_2;
  reg        [7:0]    _5_2_inner_activation;
  reg        [7:0]    _5_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_2_inner_macOut;

  assign _zz__zz__5_2_inner_macOut = ($signed(io_mulInput) * $signed(_5_2_inner_activation));
  assign _zz__zz__5_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_2_inner_macOut)) ? 16'h007f : _zz__5_2_inner_macOut_2);
  assign _zz__5_2_inner_macOut_2 = (($signed(_zz__5_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_2_inner_activation;
    end else begin
      io_macOut = _5_2_inner_macOut;
    end
  end

  assign _zz__5_2_inner_macOut = ($signed(_zz__zz__5_2_inner_macOut) + $signed(_zz__zz__5_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_2_inner_activation <= 8'h00;
      _5_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_2_inner_activation <= io_addInput;
      end else begin
        _5_2_inner_macOut <= _zz__5_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_161 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_1_inner_macOut;
  wire       [15:0]   _zz__zz__5_1_inner_macOut_1;
  wire       [15:0]   _zz__5_1_inner_macOut_1;
  wire       [15:0]   _zz__5_1_inner_macOut_2;
  reg        [7:0]    _5_1_inner_activation;
  reg        [7:0]    _5_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_1_inner_macOut;

  assign _zz__zz__5_1_inner_macOut = ($signed(io_mulInput) * $signed(_5_1_inner_activation));
  assign _zz__zz__5_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_1_inner_macOut)) ? 16'h007f : _zz__5_1_inner_macOut_2);
  assign _zz__5_1_inner_macOut_2 = (($signed(_zz__5_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_1_inner_activation;
    end else begin
      io_macOut = _5_1_inner_macOut;
    end
  end

  assign _zz__5_1_inner_macOut = ($signed(_zz__zz__5_1_inner_macOut) + $signed(_zz__zz__5_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_1_inner_activation <= 8'h00;
      _5_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_1_inner_activation <= io_addInput;
      end else begin
        _5_1_inner_macOut <= _zz__5_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_160 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__5_0_inner_macOut;
  wire       [15:0]   _zz__zz__5_0_inner_macOut_1;
  wire       [15:0]   _zz__5_0_inner_macOut_1;
  wire       [15:0]   _zz__5_0_inner_macOut_2;
  reg        [7:0]    _5_0_inner_activation;
  reg        [7:0]    _5_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__5_0_inner_macOut;

  assign _zz__zz__5_0_inner_macOut = ($signed(io_mulInput) * $signed(_5_0_inner_activation));
  assign _zz__zz__5_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__5_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__5_0_inner_macOut)) ? 16'h007f : _zz__5_0_inner_macOut_2);
  assign _zz__5_0_inner_macOut_2 = (($signed(_zz__5_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__5_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _5_0_inner_activation;
    end else begin
      io_macOut = _5_0_inner_macOut;
    end
  end

  assign _zz__5_0_inner_macOut = ($signed(_zz__zz__5_0_inner_macOut) + $signed(_zz__zz__5_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _5_0_inner_activation <= 8'h00;
      _5_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _5_0_inner_activation <= io_addInput;
      end else begin
        _5_0_inner_macOut <= _zz__5_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_159 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_31_inner_macOut;
  wire       [15:0]   _zz__zz__4_31_inner_macOut_1;
  wire       [15:0]   _zz__4_31_inner_macOut_1;
  wire       [15:0]   _zz__4_31_inner_macOut_2;
  reg        [7:0]    _4_31_inner_activation;
  reg        [7:0]    _4_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_31_inner_macOut;

  assign _zz__zz__4_31_inner_macOut = ($signed(io_mulInput) * $signed(_4_31_inner_activation));
  assign _zz__zz__4_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_31_inner_macOut)) ? 16'h007f : _zz__4_31_inner_macOut_2);
  assign _zz__4_31_inner_macOut_2 = (($signed(_zz__4_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_31_inner_activation;
    end else begin
      io_macOut = _4_31_inner_macOut;
    end
  end

  assign _zz__4_31_inner_macOut = ($signed(_zz__zz__4_31_inner_macOut) + $signed(_zz__zz__4_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_31_inner_activation <= 8'h00;
      _4_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_31_inner_activation <= io_addInput;
      end else begin
        _4_31_inner_macOut <= _zz__4_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_158 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_30_inner_macOut;
  wire       [15:0]   _zz__zz__4_30_inner_macOut_1;
  wire       [15:0]   _zz__4_30_inner_macOut_1;
  wire       [15:0]   _zz__4_30_inner_macOut_2;
  reg        [7:0]    _4_30_inner_activation;
  reg        [7:0]    _4_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_30_inner_macOut;

  assign _zz__zz__4_30_inner_macOut = ($signed(io_mulInput) * $signed(_4_30_inner_activation));
  assign _zz__zz__4_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_30_inner_macOut)) ? 16'h007f : _zz__4_30_inner_macOut_2);
  assign _zz__4_30_inner_macOut_2 = (($signed(_zz__4_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_30_inner_activation;
    end else begin
      io_macOut = _4_30_inner_macOut;
    end
  end

  assign _zz__4_30_inner_macOut = ($signed(_zz__zz__4_30_inner_macOut) + $signed(_zz__zz__4_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_30_inner_activation <= 8'h00;
      _4_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_30_inner_activation <= io_addInput;
      end else begin
        _4_30_inner_macOut <= _zz__4_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_157 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_29_inner_macOut;
  wire       [15:0]   _zz__zz__4_29_inner_macOut_1;
  wire       [15:0]   _zz__4_29_inner_macOut_1;
  wire       [15:0]   _zz__4_29_inner_macOut_2;
  reg        [7:0]    _4_29_inner_activation;
  reg        [7:0]    _4_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_29_inner_macOut;

  assign _zz__zz__4_29_inner_macOut = ($signed(io_mulInput) * $signed(_4_29_inner_activation));
  assign _zz__zz__4_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_29_inner_macOut)) ? 16'h007f : _zz__4_29_inner_macOut_2);
  assign _zz__4_29_inner_macOut_2 = (($signed(_zz__4_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_29_inner_activation;
    end else begin
      io_macOut = _4_29_inner_macOut;
    end
  end

  assign _zz__4_29_inner_macOut = ($signed(_zz__zz__4_29_inner_macOut) + $signed(_zz__zz__4_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_29_inner_activation <= 8'h00;
      _4_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_29_inner_activation <= io_addInput;
      end else begin
        _4_29_inner_macOut <= _zz__4_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_156 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_28_inner_macOut;
  wire       [15:0]   _zz__zz__4_28_inner_macOut_1;
  wire       [15:0]   _zz__4_28_inner_macOut_1;
  wire       [15:0]   _zz__4_28_inner_macOut_2;
  reg        [7:0]    _4_28_inner_activation;
  reg        [7:0]    _4_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_28_inner_macOut;

  assign _zz__zz__4_28_inner_macOut = ($signed(io_mulInput) * $signed(_4_28_inner_activation));
  assign _zz__zz__4_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_28_inner_macOut)) ? 16'h007f : _zz__4_28_inner_macOut_2);
  assign _zz__4_28_inner_macOut_2 = (($signed(_zz__4_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_28_inner_activation;
    end else begin
      io_macOut = _4_28_inner_macOut;
    end
  end

  assign _zz__4_28_inner_macOut = ($signed(_zz__zz__4_28_inner_macOut) + $signed(_zz__zz__4_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_28_inner_activation <= 8'h00;
      _4_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_28_inner_activation <= io_addInput;
      end else begin
        _4_28_inner_macOut <= _zz__4_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_155 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_27_inner_macOut;
  wire       [15:0]   _zz__zz__4_27_inner_macOut_1;
  wire       [15:0]   _zz__4_27_inner_macOut_1;
  wire       [15:0]   _zz__4_27_inner_macOut_2;
  reg        [7:0]    _4_27_inner_activation;
  reg        [7:0]    _4_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_27_inner_macOut;

  assign _zz__zz__4_27_inner_macOut = ($signed(io_mulInput) * $signed(_4_27_inner_activation));
  assign _zz__zz__4_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_27_inner_macOut)) ? 16'h007f : _zz__4_27_inner_macOut_2);
  assign _zz__4_27_inner_macOut_2 = (($signed(_zz__4_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_27_inner_activation;
    end else begin
      io_macOut = _4_27_inner_macOut;
    end
  end

  assign _zz__4_27_inner_macOut = ($signed(_zz__zz__4_27_inner_macOut) + $signed(_zz__zz__4_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_27_inner_activation <= 8'h00;
      _4_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_27_inner_activation <= io_addInput;
      end else begin
        _4_27_inner_macOut <= _zz__4_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_154 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_26_inner_macOut;
  wire       [15:0]   _zz__zz__4_26_inner_macOut_1;
  wire       [15:0]   _zz__4_26_inner_macOut_1;
  wire       [15:0]   _zz__4_26_inner_macOut_2;
  reg        [7:0]    _4_26_inner_activation;
  reg        [7:0]    _4_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_26_inner_macOut;

  assign _zz__zz__4_26_inner_macOut = ($signed(io_mulInput) * $signed(_4_26_inner_activation));
  assign _zz__zz__4_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_26_inner_macOut)) ? 16'h007f : _zz__4_26_inner_macOut_2);
  assign _zz__4_26_inner_macOut_2 = (($signed(_zz__4_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_26_inner_activation;
    end else begin
      io_macOut = _4_26_inner_macOut;
    end
  end

  assign _zz__4_26_inner_macOut = ($signed(_zz__zz__4_26_inner_macOut) + $signed(_zz__zz__4_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_26_inner_activation <= 8'h00;
      _4_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_26_inner_activation <= io_addInput;
      end else begin
        _4_26_inner_macOut <= _zz__4_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_153 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_25_inner_macOut;
  wire       [15:0]   _zz__zz__4_25_inner_macOut_1;
  wire       [15:0]   _zz__4_25_inner_macOut_1;
  wire       [15:0]   _zz__4_25_inner_macOut_2;
  reg        [7:0]    _4_25_inner_activation;
  reg        [7:0]    _4_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_25_inner_macOut;

  assign _zz__zz__4_25_inner_macOut = ($signed(io_mulInput) * $signed(_4_25_inner_activation));
  assign _zz__zz__4_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_25_inner_macOut)) ? 16'h007f : _zz__4_25_inner_macOut_2);
  assign _zz__4_25_inner_macOut_2 = (($signed(_zz__4_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_25_inner_activation;
    end else begin
      io_macOut = _4_25_inner_macOut;
    end
  end

  assign _zz__4_25_inner_macOut = ($signed(_zz__zz__4_25_inner_macOut) + $signed(_zz__zz__4_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_25_inner_activation <= 8'h00;
      _4_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_25_inner_activation <= io_addInput;
      end else begin
        _4_25_inner_macOut <= _zz__4_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_152 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_24_inner_macOut;
  wire       [15:0]   _zz__zz__4_24_inner_macOut_1;
  wire       [15:0]   _zz__4_24_inner_macOut_1;
  wire       [15:0]   _zz__4_24_inner_macOut_2;
  reg        [7:0]    _4_24_inner_activation;
  reg        [7:0]    _4_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_24_inner_macOut;

  assign _zz__zz__4_24_inner_macOut = ($signed(io_mulInput) * $signed(_4_24_inner_activation));
  assign _zz__zz__4_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_24_inner_macOut)) ? 16'h007f : _zz__4_24_inner_macOut_2);
  assign _zz__4_24_inner_macOut_2 = (($signed(_zz__4_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_24_inner_activation;
    end else begin
      io_macOut = _4_24_inner_macOut;
    end
  end

  assign _zz__4_24_inner_macOut = ($signed(_zz__zz__4_24_inner_macOut) + $signed(_zz__zz__4_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_24_inner_activation <= 8'h00;
      _4_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_24_inner_activation <= io_addInput;
      end else begin
        _4_24_inner_macOut <= _zz__4_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_151 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_23_inner_macOut;
  wire       [15:0]   _zz__zz__4_23_inner_macOut_1;
  wire       [15:0]   _zz__4_23_inner_macOut_1;
  wire       [15:0]   _zz__4_23_inner_macOut_2;
  reg        [7:0]    _4_23_inner_activation;
  reg        [7:0]    _4_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_23_inner_macOut;

  assign _zz__zz__4_23_inner_macOut = ($signed(io_mulInput) * $signed(_4_23_inner_activation));
  assign _zz__zz__4_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_23_inner_macOut)) ? 16'h007f : _zz__4_23_inner_macOut_2);
  assign _zz__4_23_inner_macOut_2 = (($signed(_zz__4_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_23_inner_activation;
    end else begin
      io_macOut = _4_23_inner_macOut;
    end
  end

  assign _zz__4_23_inner_macOut = ($signed(_zz__zz__4_23_inner_macOut) + $signed(_zz__zz__4_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_23_inner_activation <= 8'h00;
      _4_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_23_inner_activation <= io_addInput;
      end else begin
        _4_23_inner_macOut <= _zz__4_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_150 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_22_inner_macOut;
  wire       [15:0]   _zz__zz__4_22_inner_macOut_1;
  wire       [15:0]   _zz__4_22_inner_macOut_1;
  wire       [15:0]   _zz__4_22_inner_macOut_2;
  reg        [7:0]    _4_22_inner_activation;
  reg        [7:0]    _4_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_22_inner_macOut;

  assign _zz__zz__4_22_inner_macOut = ($signed(io_mulInput) * $signed(_4_22_inner_activation));
  assign _zz__zz__4_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_22_inner_macOut)) ? 16'h007f : _zz__4_22_inner_macOut_2);
  assign _zz__4_22_inner_macOut_2 = (($signed(_zz__4_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_22_inner_activation;
    end else begin
      io_macOut = _4_22_inner_macOut;
    end
  end

  assign _zz__4_22_inner_macOut = ($signed(_zz__zz__4_22_inner_macOut) + $signed(_zz__zz__4_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_22_inner_activation <= 8'h00;
      _4_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_22_inner_activation <= io_addInput;
      end else begin
        _4_22_inner_macOut <= _zz__4_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_149 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_21_inner_macOut;
  wire       [15:0]   _zz__zz__4_21_inner_macOut_1;
  wire       [15:0]   _zz__4_21_inner_macOut_1;
  wire       [15:0]   _zz__4_21_inner_macOut_2;
  reg        [7:0]    _4_21_inner_activation;
  reg        [7:0]    _4_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_21_inner_macOut;

  assign _zz__zz__4_21_inner_macOut = ($signed(io_mulInput) * $signed(_4_21_inner_activation));
  assign _zz__zz__4_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_21_inner_macOut)) ? 16'h007f : _zz__4_21_inner_macOut_2);
  assign _zz__4_21_inner_macOut_2 = (($signed(_zz__4_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_21_inner_activation;
    end else begin
      io_macOut = _4_21_inner_macOut;
    end
  end

  assign _zz__4_21_inner_macOut = ($signed(_zz__zz__4_21_inner_macOut) + $signed(_zz__zz__4_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_21_inner_activation <= 8'h00;
      _4_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_21_inner_activation <= io_addInput;
      end else begin
        _4_21_inner_macOut <= _zz__4_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_148 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_20_inner_macOut;
  wire       [15:0]   _zz__zz__4_20_inner_macOut_1;
  wire       [15:0]   _zz__4_20_inner_macOut_1;
  wire       [15:0]   _zz__4_20_inner_macOut_2;
  reg        [7:0]    _4_20_inner_activation;
  reg        [7:0]    _4_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_20_inner_macOut;

  assign _zz__zz__4_20_inner_macOut = ($signed(io_mulInput) * $signed(_4_20_inner_activation));
  assign _zz__zz__4_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_20_inner_macOut)) ? 16'h007f : _zz__4_20_inner_macOut_2);
  assign _zz__4_20_inner_macOut_2 = (($signed(_zz__4_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_20_inner_activation;
    end else begin
      io_macOut = _4_20_inner_macOut;
    end
  end

  assign _zz__4_20_inner_macOut = ($signed(_zz__zz__4_20_inner_macOut) + $signed(_zz__zz__4_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_20_inner_activation <= 8'h00;
      _4_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_20_inner_activation <= io_addInput;
      end else begin
        _4_20_inner_macOut <= _zz__4_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_147 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_19_inner_macOut;
  wire       [15:0]   _zz__zz__4_19_inner_macOut_1;
  wire       [15:0]   _zz__4_19_inner_macOut_1;
  wire       [15:0]   _zz__4_19_inner_macOut_2;
  reg        [7:0]    _4_19_inner_activation;
  reg        [7:0]    _4_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_19_inner_macOut;

  assign _zz__zz__4_19_inner_macOut = ($signed(io_mulInput) * $signed(_4_19_inner_activation));
  assign _zz__zz__4_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_19_inner_macOut)) ? 16'h007f : _zz__4_19_inner_macOut_2);
  assign _zz__4_19_inner_macOut_2 = (($signed(_zz__4_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_19_inner_activation;
    end else begin
      io_macOut = _4_19_inner_macOut;
    end
  end

  assign _zz__4_19_inner_macOut = ($signed(_zz__zz__4_19_inner_macOut) + $signed(_zz__zz__4_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_19_inner_activation <= 8'h00;
      _4_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_19_inner_activation <= io_addInput;
      end else begin
        _4_19_inner_macOut <= _zz__4_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_146 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_18_inner_macOut;
  wire       [15:0]   _zz__zz__4_18_inner_macOut_1;
  wire       [15:0]   _zz__4_18_inner_macOut_1;
  wire       [15:0]   _zz__4_18_inner_macOut_2;
  reg        [7:0]    _4_18_inner_activation;
  reg        [7:0]    _4_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_18_inner_macOut;

  assign _zz__zz__4_18_inner_macOut = ($signed(io_mulInput) * $signed(_4_18_inner_activation));
  assign _zz__zz__4_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_18_inner_macOut)) ? 16'h007f : _zz__4_18_inner_macOut_2);
  assign _zz__4_18_inner_macOut_2 = (($signed(_zz__4_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_18_inner_activation;
    end else begin
      io_macOut = _4_18_inner_macOut;
    end
  end

  assign _zz__4_18_inner_macOut = ($signed(_zz__zz__4_18_inner_macOut) + $signed(_zz__zz__4_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_18_inner_activation <= 8'h00;
      _4_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_18_inner_activation <= io_addInput;
      end else begin
        _4_18_inner_macOut <= _zz__4_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_145 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_17_inner_macOut;
  wire       [15:0]   _zz__zz__4_17_inner_macOut_1;
  wire       [15:0]   _zz__4_17_inner_macOut_1;
  wire       [15:0]   _zz__4_17_inner_macOut_2;
  reg        [7:0]    _4_17_inner_activation;
  reg        [7:0]    _4_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_17_inner_macOut;

  assign _zz__zz__4_17_inner_macOut = ($signed(io_mulInput) * $signed(_4_17_inner_activation));
  assign _zz__zz__4_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_17_inner_macOut)) ? 16'h007f : _zz__4_17_inner_macOut_2);
  assign _zz__4_17_inner_macOut_2 = (($signed(_zz__4_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_17_inner_activation;
    end else begin
      io_macOut = _4_17_inner_macOut;
    end
  end

  assign _zz__4_17_inner_macOut = ($signed(_zz__zz__4_17_inner_macOut) + $signed(_zz__zz__4_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_17_inner_activation <= 8'h00;
      _4_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_17_inner_activation <= io_addInput;
      end else begin
        _4_17_inner_macOut <= _zz__4_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_144 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_16_inner_macOut;
  wire       [15:0]   _zz__zz__4_16_inner_macOut_1;
  wire       [15:0]   _zz__4_16_inner_macOut_1;
  wire       [15:0]   _zz__4_16_inner_macOut_2;
  reg        [7:0]    _4_16_inner_activation;
  reg        [7:0]    _4_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_16_inner_macOut;

  assign _zz__zz__4_16_inner_macOut = ($signed(io_mulInput) * $signed(_4_16_inner_activation));
  assign _zz__zz__4_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_16_inner_macOut)) ? 16'h007f : _zz__4_16_inner_macOut_2);
  assign _zz__4_16_inner_macOut_2 = (($signed(_zz__4_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_16_inner_activation;
    end else begin
      io_macOut = _4_16_inner_macOut;
    end
  end

  assign _zz__4_16_inner_macOut = ($signed(_zz__zz__4_16_inner_macOut) + $signed(_zz__zz__4_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_16_inner_activation <= 8'h00;
      _4_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_16_inner_activation <= io_addInput;
      end else begin
        _4_16_inner_macOut <= _zz__4_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_143 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_15_inner_macOut;
  wire       [15:0]   _zz__zz__4_15_inner_macOut_1;
  wire       [15:0]   _zz__4_15_inner_macOut_1;
  wire       [15:0]   _zz__4_15_inner_macOut_2;
  reg        [7:0]    _4_15_inner_activation;
  reg        [7:0]    _4_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_15_inner_macOut;

  assign _zz__zz__4_15_inner_macOut = ($signed(io_mulInput) * $signed(_4_15_inner_activation));
  assign _zz__zz__4_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_15_inner_macOut)) ? 16'h007f : _zz__4_15_inner_macOut_2);
  assign _zz__4_15_inner_macOut_2 = (($signed(_zz__4_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_15_inner_activation;
    end else begin
      io_macOut = _4_15_inner_macOut;
    end
  end

  assign _zz__4_15_inner_macOut = ($signed(_zz__zz__4_15_inner_macOut) + $signed(_zz__zz__4_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_15_inner_activation <= 8'h00;
      _4_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_15_inner_activation <= io_addInput;
      end else begin
        _4_15_inner_macOut <= _zz__4_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_142 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_14_inner_macOut;
  wire       [15:0]   _zz__zz__4_14_inner_macOut_1;
  wire       [15:0]   _zz__4_14_inner_macOut_1;
  wire       [15:0]   _zz__4_14_inner_macOut_2;
  reg        [7:0]    _4_14_inner_activation;
  reg        [7:0]    _4_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_14_inner_macOut;

  assign _zz__zz__4_14_inner_macOut = ($signed(io_mulInput) * $signed(_4_14_inner_activation));
  assign _zz__zz__4_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_14_inner_macOut)) ? 16'h007f : _zz__4_14_inner_macOut_2);
  assign _zz__4_14_inner_macOut_2 = (($signed(_zz__4_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_14_inner_activation;
    end else begin
      io_macOut = _4_14_inner_macOut;
    end
  end

  assign _zz__4_14_inner_macOut = ($signed(_zz__zz__4_14_inner_macOut) + $signed(_zz__zz__4_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_14_inner_activation <= 8'h00;
      _4_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_14_inner_activation <= io_addInput;
      end else begin
        _4_14_inner_macOut <= _zz__4_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_141 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_13_inner_macOut;
  wire       [15:0]   _zz__zz__4_13_inner_macOut_1;
  wire       [15:0]   _zz__4_13_inner_macOut_1;
  wire       [15:0]   _zz__4_13_inner_macOut_2;
  reg        [7:0]    _4_13_inner_activation;
  reg        [7:0]    _4_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_13_inner_macOut;

  assign _zz__zz__4_13_inner_macOut = ($signed(io_mulInput) * $signed(_4_13_inner_activation));
  assign _zz__zz__4_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_13_inner_macOut)) ? 16'h007f : _zz__4_13_inner_macOut_2);
  assign _zz__4_13_inner_macOut_2 = (($signed(_zz__4_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_13_inner_activation;
    end else begin
      io_macOut = _4_13_inner_macOut;
    end
  end

  assign _zz__4_13_inner_macOut = ($signed(_zz__zz__4_13_inner_macOut) + $signed(_zz__zz__4_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_13_inner_activation <= 8'h00;
      _4_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_13_inner_activation <= io_addInput;
      end else begin
        _4_13_inner_macOut <= _zz__4_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_140 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_12_inner_macOut;
  wire       [15:0]   _zz__zz__4_12_inner_macOut_1;
  wire       [15:0]   _zz__4_12_inner_macOut_1;
  wire       [15:0]   _zz__4_12_inner_macOut_2;
  reg        [7:0]    _4_12_inner_activation;
  reg        [7:0]    _4_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_12_inner_macOut;

  assign _zz__zz__4_12_inner_macOut = ($signed(io_mulInput) * $signed(_4_12_inner_activation));
  assign _zz__zz__4_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_12_inner_macOut)) ? 16'h007f : _zz__4_12_inner_macOut_2);
  assign _zz__4_12_inner_macOut_2 = (($signed(_zz__4_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_12_inner_activation;
    end else begin
      io_macOut = _4_12_inner_macOut;
    end
  end

  assign _zz__4_12_inner_macOut = ($signed(_zz__zz__4_12_inner_macOut) + $signed(_zz__zz__4_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_12_inner_activation <= 8'h00;
      _4_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_12_inner_activation <= io_addInput;
      end else begin
        _4_12_inner_macOut <= _zz__4_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_139 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_11_inner_macOut;
  wire       [15:0]   _zz__zz__4_11_inner_macOut_1;
  wire       [15:0]   _zz__4_11_inner_macOut_1;
  wire       [15:0]   _zz__4_11_inner_macOut_2;
  reg        [7:0]    _4_11_inner_activation;
  reg        [7:0]    _4_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_11_inner_macOut;

  assign _zz__zz__4_11_inner_macOut = ($signed(io_mulInput) * $signed(_4_11_inner_activation));
  assign _zz__zz__4_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_11_inner_macOut)) ? 16'h007f : _zz__4_11_inner_macOut_2);
  assign _zz__4_11_inner_macOut_2 = (($signed(_zz__4_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_11_inner_activation;
    end else begin
      io_macOut = _4_11_inner_macOut;
    end
  end

  assign _zz__4_11_inner_macOut = ($signed(_zz__zz__4_11_inner_macOut) + $signed(_zz__zz__4_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_11_inner_activation <= 8'h00;
      _4_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_11_inner_activation <= io_addInput;
      end else begin
        _4_11_inner_macOut <= _zz__4_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_138 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_10_inner_macOut;
  wire       [15:0]   _zz__zz__4_10_inner_macOut_1;
  wire       [15:0]   _zz__4_10_inner_macOut_1;
  wire       [15:0]   _zz__4_10_inner_macOut_2;
  reg        [7:0]    _4_10_inner_activation;
  reg        [7:0]    _4_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_10_inner_macOut;

  assign _zz__zz__4_10_inner_macOut = ($signed(io_mulInput) * $signed(_4_10_inner_activation));
  assign _zz__zz__4_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_10_inner_macOut)) ? 16'h007f : _zz__4_10_inner_macOut_2);
  assign _zz__4_10_inner_macOut_2 = (($signed(_zz__4_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_10_inner_activation;
    end else begin
      io_macOut = _4_10_inner_macOut;
    end
  end

  assign _zz__4_10_inner_macOut = ($signed(_zz__zz__4_10_inner_macOut) + $signed(_zz__zz__4_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_10_inner_activation <= 8'h00;
      _4_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_10_inner_activation <= io_addInput;
      end else begin
        _4_10_inner_macOut <= _zz__4_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_137 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_9_inner_macOut;
  wire       [15:0]   _zz__zz__4_9_inner_macOut_1;
  wire       [15:0]   _zz__4_9_inner_macOut_1;
  wire       [15:0]   _zz__4_9_inner_macOut_2;
  reg        [7:0]    _4_9_inner_activation;
  reg        [7:0]    _4_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_9_inner_macOut;

  assign _zz__zz__4_9_inner_macOut = ($signed(io_mulInput) * $signed(_4_9_inner_activation));
  assign _zz__zz__4_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_9_inner_macOut)) ? 16'h007f : _zz__4_9_inner_macOut_2);
  assign _zz__4_9_inner_macOut_2 = (($signed(_zz__4_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_9_inner_activation;
    end else begin
      io_macOut = _4_9_inner_macOut;
    end
  end

  assign _zz__4_9_inner_macOut = ($signed(_zz__zz__4_9_inner_macOut) + $signed(_zz__zz__4_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_9_inner_activation <= 8'h00;
      _4_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_9_inner_activation <= io_addInput;
      end else begin
        _4_9_inner_macOut <= _zz__4_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_136 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_8_inner_macOut;
  wire       [15:0]   _zz__zz__4_8_inner_macOut_1;
  wire       [15:0]   _zz__4_8_inner_macOut_1;
  wire       [15:0]   _zz__4_8_inner_macOut_2;
  reg        [7:0]    _4_8_inner_activation;
  reg        [7:0]    _4_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_8_inner_macOut;

  assign _zz__zz__4_8_inner_macOut = ($signed(io_mulInput) * $signed(_4_8_inner_activation));
  assign _zz__zz__4_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_8_inner_macOut)) ? 16'h007f : _zz__4_8_inner_macOut_2);
  assign _zz__4_8_inner_macOut_2 = (($signed(_zz__4_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_8_inner_activation;
    end else begin
      io_macOut = _4_8_inner_macOut;
    end
  end

  assign _zz__4_8_inner_macOut = ($signed(_zz__zz__4_8_inner_macOut) + $signed(_zz__zz__4_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_8_inner_activation <= 8'h00;
      _4_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_8_inner_activation <= io_addInput;
      end else begin
        _4_8_inner_macOut <= _zz__4_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_135 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_7_inner_macOut;
  wire       [15:0]   _zz__zz__4_7_inner_macOut_1;
  wire       [15:0]   _zz__4_7_inner_macOut_1;
  wire       [15:0]   _zz__4_7_inner_macOut_2;
  reg        [7:0]    _4_7_inner_activation;
  reg        [7:0]    _4_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_7_inner_macOut;

  assign _zz__zz__4_7_inner_macOut = ($signed(io_mulInput) * $signed(_4_7_inner_activation));
  assign _zz__zz__4_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_7_inner_macOut)) ? 16'h007f : _zz__4_7_inner_macOut_2);
  assign _zz__4_7_inner_macOut_2 = (($signed(_zz__4_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_7_inner_activation;
    end else begin
      io_macOut = _4_7_inner_macOut;
    end
  end

  assign _zz__4_7_inner_macOut = ($signed(_zz__zz__4_7_inner_macOut) + $signed(_zz__zz__4_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_7_inner_activation <= 8'h00;
      _4_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_7_inner_activation <= io_addInput;
      end else begin
        _4_7_inner_macOut <= _zz__4_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_134 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_6_inner_macOut;
  wire       [15:0]   _zz__zz__4_6_inner_macOut_1;
  wire       [15:0]   _zz__4_6_inner_macOut_1;
  wire       [15:0]   _zz__4_6_inner_macOut_2;
  reg        [7:0]    _4_6_inner_activation;
  reg        [7:0]    _4_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_6_inner_macOut;

  assign _zz__zz__4_6_inner_macOut = ($signed(io_mulInput) * $signed(_4_6_inner_activation));
  assign _zz__zz__4_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_6_inner_macOut)) ? 16'h007f : _zz__4_6_inner_macOut_2);
  assign _zz__4_6_inner_macOut_2 = (($signed(_zz__4_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_6_inner_activation;
    end else begin
      io_macOut = _4_6_inner_macOut;
    end
  end

  assign _zz__4_6_inner_macOut = ($signed(_zz__zz__4_6_inner_macOut) + $signed(_zz__zz__4_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_6_inner_activation <= 8'h00;
      _4_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_6_inner_activation <= io_addInput;
      end else begin
        _4_6_inner_macOut <= _zz__4_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_133 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_5_inner_macOut;
  wire       [15:0]   _zz__zz__4_5_inner_macOut_1;
  wire       [15:0]   _zz__4_5_inner_macOut_1;
  wire       [15:0]   _zz__4_5_inner_macOut_2;
  reg        [7:0]    _4_5_inner_activation;
  reg        [7:0]    _4_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_5_inner_macOut;

  assign _zz__zz__4_5_inner_macOut = ($signed(io_mulInput) * $signed(_4_5_inner_activation));
  assign _zz__zz__4_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_5_inner_macOut)) ? 16'h007f : _zz__4_5_inner_macOut_2);
  assign _zz__4_5_inner_macOut_2 = (($signed(_zz__4_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_5_inner_activation;
    end else begin
      io_macOut = _4_5_inner_macOut;
    end
  end

  assign _zz__4_5_inner_macOut = ($signed(_zz__zz__4_5_inner_macOut) + $signed(_zz__zz__4_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_5_inner_activation <= 8'h00;
      _4_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_5_inner_activation <= io_addInput;
      end else begin
        _4_5_inner_macOut <= _zz__4_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_132 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_4_inner_macOut;
  wire       [15:0]   _zz__zz__4_4_inner_macOut_1;
  wire       [15:0]   _zz__4_4_inner_macOut_1;
  wire       [15:0]   _zz__4_4_inner_macOut_2;
  reg        [7:0]    _4_4_inner_activation;
  reg        [7:0]    _4_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_4_inner_macOut;

  assign _zz__zz__4_4_inner_macOut = ($signed(io_mulInput) * $signed(_4_4_inner_activation));
  assign _zz__zz__4_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_4_inner_macOut)) ? 16'h007f : _zz__4_4_inner_macOut_2);
  assign _zz__4_4_inner_macOut_2 = (($signed(_zz__4_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_4_inner_activation;
    end else begin
      io_macOut = _4_4_inner_macOut;
    end
  end

  assign _zz__4_4_inner_macOut = ($signed(_zz__zz__4_4_inner_macOut) + $signed(_zz__zz__4_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_4_inner_activation <= 8'h00;
      _4_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_4_inner_activation <= io_addInput;
      end else begin
        _4_4_inner_macOut <= _zz__4_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_131 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_3_inner_macOut;
  wire       [15:0]   _zz__zz__4_3_inner_macOut_1;
  wire       [15:0]   _zz__4_3_inner_macOut_1;
  wire       [15:0]   _zz__4_3_inner_macOut_2;
  reg        [7:0]    _4_3_inner_activation;
  reg        [7:0]    _4_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_3_inner_macOut;

  assign _zz__zz__4_3_inner_macOut = ($signed(io_mulInput) * $signed(_4_3_inner_activation));
  assign _zz__zz__4_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_3_inner_macOut)) ? 16'h007f : _zz__4_3_inner_macOut_2);
  assign _zz__4_3_inner_macOut_2 = (($signed(_zz__4_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_3_inner_activation;
    end else begin
      io_macOut = _4_3_inner_macOut;
    end
  end

  assign _zz__4_3_inner_macOut = ($signed(_zz__zz__4_3_inner_macOut) + $signed(_zz__zz__4_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_3_inner_activation <= 8'h00;
      _4_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_3_inner_activation <= io_addInput;
      end else begin
        _4_3_inner_macOut <= _zz__4_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_130 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_2_inner_macOut;
  wire       [15:0]   _zz__zz__4_2_inner_macOut_1;
  wire       [15:0]   _zz__4_2_inner_macOut_1;
  wire       [15:0]   _zz__4_2_inner_macOut_2;
  reg        [7:0]    _4_2_inner_activation;
  reg        [7:0]    _4_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_2_inner_macOut;

  assign _zz__zz__4_2_inner_macOut = ($signed(io_mulInput) * $signed(_4_2_inner_activation));
  assign _zz__zz__4_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_2_inner_macOut)) ? 16'h007f : _zz__4_2_inner_macOut_2);
  assign _zz__4_2_inner_macOut_2 = (($signed(_zz__4_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_2_inner_activation;
    end else begin
      io_macOut = _4_2_inner_macOut;
    end
  end

  assign _zz__4_2_inner_macOut = ($signed(_zz__zz__4_2_inner_macOut) + $signed(_zz__zz__4_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_2_inner_activation <= 8'h00;
      _4_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_2_inner_activation <= io_addInput;
      end else begin
        _4_2_inner_macOut <= _zz__4_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_129 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_1_inner_macOut;
  wire       [15:0]   _zz__zz__4_1_inner_macOut_1;
  wire       [15:0]   _zz__4_1_inner_macOut_1;
  wire       [15:0]   _zz__4_1_inner_macOut_2;
  reg        [7:0]    _4_1_inner_activation;
  reg        [7:0]    _4_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_1_inner_macOut;

  assign _zz__zz__4_1_inner_macOut = ($signed(io_mulInput) * $signed(_4_1_inner_activation));
  assign _zz__zz__4_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_1_inner_macOut)) ? 16'h007f : _zz__4_1_inner_macOut_2);
  assign _zz__4_1_inner_macOut_2 = (($signed(_zz__4_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_1_inner_activation;
    end else begin
      io_macOut = _4_1_inner_macOut;
    end
  end

  assign _zz__4_1_inner_macOut = ($signed(_zz__zz__4_1_inner_macOut) + $signed(_zz__zz__4_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_1_inner_activation <= 8'h00;
      _4_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_1_inner_activation <= io_addInput;
      end else begin
        _4_1_inner_macOut <= _zz__4_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_128 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__4_0_inner_macOut;
  wire       [15:0]   _zz__zz__4_0_inner_macOut_1;
  wire       [15:0]   _zz__4_0_inner_macOut_1;
  wire       [15:0]   _zz__4_0_inner_macOut_2;
  reg        [7:0]    _4_0_inner_activation;
  reg        [7:0]    _4_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__4_0_inner_macOut;

  assign _zz__zz__4_0_inner_macOut = ($signed(io_mulInput) * $signed(_4_0_inner_activation));
  assign _zz__zz__4_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__4_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__4_0_inner_macOut)) ? 16'h007f : _zz__4_0_inner_macOut_2);
  assign _zz__4_0_inner_macOut_2 = (($signed(_zz__4_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__4_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _4_0_inner_activation;
    end else begin
      io_macOut = _4_0_inner_macOut;
    end
  end

  assign _zz__4_0_inner_macOut = ($signed(_zz__zz__4_0_inner_macOut) + $signed(_zz__zz__4_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _4_0_inner_activation <= 8'h00;
      _4_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _4_0_inner_activation <= io_addInput;
      end else begin
        _4_0_inner_macOut <= _zz__4_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_127 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_31_inner_macOut;
  wire       [15:0]   _zz__zz__3_31_inner_macOut_1;
  wire       [15:0]   _zz__3_31_inner_macOut_1;
  wire       [15:0]   _zz__3_31_inner_macOut_2;
  reg        [7:0]    _3_31_inner_activation;
  reg        [7:0]    _3_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_31_inner_macOut;

  assign _zz__zz__3_31_inner_macOut = ($signed(io_mulInput) * $signed(_3_31_inner_activation));
  assign _zz__zz__3_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_31_inner_macOut)) ? 16'h007f : _zz__3_31_inner_macOut_2);
  assign _zz__3_31_inner_macOut_2 = (($signed(_zz__3_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_31_inner_activation;
    end else begin
      io_macOut = _3_31_inner_macOut;
    end
  end

  assign _zz__3_31_inner_macOut = ($signed(_zz__zz__3_31_inner_macOut) + $signed(_zz__zz__3_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_31_inner_activation <= 8'h00;
      _3_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_31_inner_activation <= io_addInput;
      end else begin
        _3_31_inner_macOut <= _zz__3_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_126 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_30_inner_macOut;
  wire       [15:0]   _zz__zz__3_30_inner_macOut_1;
  wire       [15:0]   _zz__3_30_inner_macOut_1;
  wire       [15:0]   _zz__3_30_inner_macOut_2;
  reg        [7:0]    _3_30_inner_activation;
  reg        [7:0]    _3_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_30_inner_macOut;

  assign _zz__zz__3_30_inner_macOut = ($signed(io_mulInput) * $signed(_3_30_inner_activation));
  assign _zz__zz__3_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_30_inner_macOut)) ? 16'h007f : _zz__3_30_inner_macOut_2);
  assign _zz__3_30_inner_macOut_2 = (($signed(_zz__3_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_30_inner_activation;
    end else begin
      io_macOut = _3_30_inner_macOut;
    end
  end

  assign _zz__3_30_inner_macOut = ($signed(_zz__zz__3_30_inner_macOut) + $signed(_zz__zz__3_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_30_inner_activation <= 8'h00;
      _3_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_30_inner_activation <= io_addInput;
      end else begin
        _3_30_inner_macOut <= _zz__3_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_125 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_29_inner_macOut;
  wire       [15:0]   _zz__zz__3_29_inner_macOut_1;
  wire       [15:0]   _zz__3_29_inner_macOut_1;
  wire       [15:0]   _zz__3_29_inner_macOut_2;
  reg        [7:0]    _3_29_inner_activation;
  reg        [7:0]    _3_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_29_inner_macOut;

  assign _zz__zz__3_29_inner_macOut = ($signed(io_mulInput) * $signed(_3_29_inner_activation));
  assign _zz__zz__3_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_29_inner_macOut)) ? 16'h007f : _zz__3_29_inner_macOut_2);
  assign _zz__3_29_inner_macOut_2 = (($signed(_zz__3_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_29_inner_activation;
    end else begin
      io_macOut = _3_29_inner_macOut;
    end
  end

  assign _zz__3_29_inner_macOut = ($signed(_zz__zz__3_29_inner_macOut) + $signed(_zz__zz__3_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_29_inner_activation <= 8'h00;
      _3_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_29_inner_activation <= io_addInput;
      end else begin
        _3_29_inner_macOut <= _zz__3_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_124 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_28_inner_macOut;
  wire       [15:0]   _zz__zz__3_28_inner_macOut_1;
  wire       [15:0]   _zz__3_28_inner_macOut_1;
  wire       [15:0]   _zz__3_28_inner_macOut_2;
  reg        [7:0]    _3_28_inner_activation;
  reg        [7:0]    _3_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_28_inner_macOut;

  assign _zz__zz__3_28_inner_macOut = ($signed(io_mulInput) * $signed(_3_28_inner_activation));
  assign _zz__zz__3_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_28_inner_macOut)) ? 16'h007f : _zz__3_28_inner_macOut_2);
  assign _zz__3_28_inner_macOut_2 = (($signed(_zz__3_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_28_inner_activation;
    end else begin
      io_macOut = _3_28_inner_macOut;
    end
  end

  assign _zz__3_28_inner_macOut = ($signed(_zz__zz__3_28_inner_macOut) + $signed(_zz__zz__3_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_28_inner_activation <= 8'h00;
      _3_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_28_inner_activation <= io_addInput;
      end else begin
        _3_28_inner_macOut <= _zz__3_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_123 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_27_inner_macOut;
  wire       [15:0]   _zz__zz__3_27_inner_macOut_1;
  wire       [15:0]   _zz__3_27_inner_macOut_1;
  wire       [15:0]   _zz__3_27_inner_macOut_2;
  reg        [7:0]    _3_27_inner_activation;
  reg        [7:0]    _3_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_27_inner_macOut;

  assign _zz__zz__3_27_inner_macOut = ($signed(io_mulInput) * $signed(_3_27_inner_activation));
  assign _zz__zz__3_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_27_inner_macOut)) ? 16'h007f : _zz__3_27_inner_macOut_2);
  assign _zz__3_27_inner_macOut_2 = (($signed(_zz__3_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_27_inner_activation;
    end else begin
      io_macOut = _3_27_inner_macOut;
    end
  end

  assign _zz__3_27_inner_macOut = ($signed(_zz__zz__3_27_inner_macOut) + $signed(_zz__zz__3_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_27_inner_activation <= 8'h00;
      _3_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_27_inner_activation <= io_addInput;
      end else begin
        _3_27_inner_macOut <= _zz__3_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_122 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_26_inner_macOut;
  wire       [15:0]   _zz__zz__3_26_inner_macOut_1;
  wire       [15:0]   _zz__3_26_inner_macOut_1;
  wire       [15:0]   _zz__3_26_inner_macOut_2;
  reg        [7:0]    _3_26_inner_activation;
  reg        [7:0]    _3_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_26_inner_macOut;

  assign _zz__zz__3_26_inner_macOut = ($signed(io_mulInput) * $signed(_3_26_inner_activation));
  assign _zz__zz__3_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_26_inner_macOut)) ? 16'h007f : _zz__3_26_inner_macOut_2);
  assign _zz__3_26_inner_macOut_2 = (($signed(_zz__3_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_26_inner_activation;
    end else begin
      io_macOut = _3_26_inner_macOut;
    end
  end

  assign _zz__3_26_inner_macOut = ($signed(_zz__zz__3_26_inner_macOut) + $signed(_zz__zz__3_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_26_inner_activation <= 8'h00;
      _3_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_26_inner_activation <= io_addInput;
      end else begin
        _3_26_inner_macOut <= _zz__3_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_121 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_25_inner_macOut;
  wire       [15:0]   _zz__zz__3_25_inner_macOut_1;
  wire       [15:0]   _zz__3_25_inner_macOut_1;
  wire       [15:0]   _zz__3_25_inner_macOut_2;
  reg        [7:0]    _3_25_inner_activation;
  reg        [7:0]    _3_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_25_inner_macOut;

  assign _zz__zz__3_25_inner_macOut = ($signed(io_mulInput) * $signed(_3_25_inner_activation));
  assign _zz__zz__3_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_25_inner_macOut)) ? 16'h007f : _zz__3_25_inner_macOut_2);
  assign _zz__3_25_inner_macOut_2 = (($signed(_zz__3_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_25_inner_activation;
    end else begin
      io_macOut = _3_25_inner_macOut;
    end
  end

  assign _zz__3_25_inner_macOut = ($signed(_zz__zz__3_25_inner_macOut) + $signed(_zz__zz__3_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_25_inner_activation <= 8'h00;
      _3_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_25_inner_activation <= io_addInput;
      end else begin
        _3_25_inner_macOut <= _zz__3_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_120 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_24_inner_macOut;
  wire       [15:0]   _zz__zz__3_24_inner_macOut_1;
  wire       [15:0]   _zz__3_24_inner_macOut_1;
  wire       [15:0]   _zz__3_24_inner_macOut_2;
  reg        [7:0]    _3_24_inner_activation;
  reg        [7:0]    _3_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_24_inner_macOut;

  assign _zz__zz__3_24_inner_macOut = ($signed(io_mulInput) * $signed(_3_24_inner_activation));
  assign _zz__zz__3_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_24_inner_macOut)) ? 16'h007f : _zz__3_24_inner_macOut_2);
  assign _zz__3_24_inner_macOut_2 = (($signed(_zz__3_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_24_inner_activation;
    end else begin
      io_macOut = _3_24_inner_macOut;
    end
  end

  assign _zz__3_24_inner_macOut = ($signed(_zz__zz__3_24_inner_macOut) + $signed(_zz__zz__3_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_24_inner_activation <= 8'h00;
      _3_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_24_inner_activation <= io_addInput;
      end else begin
        _3_24_inner_macOut <= _zz__3_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_119 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_23_inner_macOut;
  wire       [15:0]   _zz__zz__3_23_inner_macOut_1;
  wire       [15:0]   _zz__3_23_inner_macOut_1;
  wire       [15:0]   _zz__3_23_inner_macOut_2;
  reg        [7:0]    _3_23_inner_activation;
  reg        [7:0]    _3_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_23_inner_macOut;

  assign _zz__zz__3_23_inner_macOut = ($signed(io_mulInput) * $signed(_3_23_inner_activation));
  assign _zz__zz__3_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_23_inner_macOut)) ? 16'h007f : _zz__3_23_inner_macOut_2);
  assign _zz__3_23_inner_macOut_2 = (($signed(_zz__3_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_23_inner_activation;
    end else begin
      io_macOut = _3_23_inner_macOut;
    end
  end

  assign _zz__3_23_inner_macOut = ($signed(_zz__zz__3_23_inner_macOut) + $signed(_zz__zz__3_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_23_inner_activation <= 8'h00;
      _3_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_23_inner_activation <= io_addInput;
      end else begin
        _3_23_inner_macOut <= _zz__3_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_118 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_22_inner_macOut;
  wire       [15:0]   _zz__zz__3_22_inner_macOut_1;
  wire       [15:0]   _zz__3_22_inner_macOut_1;
  wire       [15:0]   _zz__3_22_inner_macOut_2;
  reg        [7:0]    _3_22_inner_activation;
  reg        [7:0]    _3_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_22_inner_macOut;

  assign _zz__zz__3_22_inner_macOut = ($signed(io_mulInput) * $signed(_3_22_inner_activation));
  assign _zz__zz__3_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_22_inner_macOut)) ? 16'h007f : _zz__3_22_inner_macOut_2);
  assign _zz__3_22_inner_macOut_2 = (($signed(_zz__3_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_22_inner_activation;
    end else begin
      io_macOut = _3_22_inner_macOut;
    end
  end

  assign _zz__3_22_inner_macOut = ($signed(_zz__zz__3_22_inner_macOut) + $signed(_zz__zz__3_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_22_inner_activation <= 8'h00;
      _3_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_22_inner_activation <= io_addInput;
      end else begin
        _3_22_inner_macOut <= _zz__3_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_117 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_21_inner_macOut;
  wire       [15:0]   _zz__zz__3_21_inner_macOut_1;
  wire       [15:0]   _zz__3_21_inner_macOut_1;
  wire       [15:0]   _zz__3_21_inner_macOut_2;
  reg        [7:0]    _3_21_inner_activation;
  reg        [7:0]    _3_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_21_inner_macOut;

  assign _zz__zz__3_21_inner_macOut = ($signed(io_mulInput) * $signed(_3_21_inner_activation));
  assign _zz__zz__3_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_21_inner_macOut)) ? 16'h007f : _zz__3_21_inner_macOut_2);
  assign _zz__3_21_inner_macOut_2 = (($signed(_zz__3_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_21_inner_activation;
    end else begin
      io_macOut = _3_21_inner_macOut;
    end
  end

  assign _zz__3_21_inner_macOut = ($signed(_zz__zz__3_21_inner_macOut) + $signed(_zz__zz__3_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_21_inner_activation <= 8'h00;
      _3_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_21_inner_activation <= io_addInput;
      end else begin
        _3_21_inner_macOut <= _zz__3_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_116 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_20_inner_macOut;
  wire       [15:0]   _zz__zz__3_20_inner_macOut_1;
  wire       [15:0]   _zz__3_20_inner_macOut_1;
  wire       [15:0]   _zz__3_20_inner_macOut_2;
  reg        [7:0]    _3_20_inner_activation;
  reg        [7:0]    _3_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_20_inner_macOut;

  assign _zz__zz__3_20_inner_macOut = ($signed(io_mulInput) * $signed(_3_20_inner_activation));
  assign _zz__zz__3_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_20_inner_macOut)) ? 16'h007f : _zz__3_20_inner_macOut_2);
  assign _zz__3_20_inner_macOut_2 = (($signed(_zz__3_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_20_inner_activation;
    end else begin
      io_macOut = _3_20_inner_macOut;
    end
  end

  assign _zz__3_20_inner_macOut = ($signed(_zz__zz__3_20_inner_macOut) + $signed(_zz__zz__3_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_20_inner_activation <= 8'h00;
      _3_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_20_inner_activation <= io_addInput;
      end else begin
        _3_20_inner_macOut <= _zz__3_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_115 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_19_inner_macOut;
  wire       [15:0]   _zz__zz__3_19_inner_macOut_1;
  wire       [15:0]   _zz__3_19_inner_macOut_1;
  wire       [15:0]   _zz__3_19_inner_macOut_2;
  reg        [7:0]    _3_19_inner_activation;
  reg        [7:0]    _3_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_19_inner_macOut;

  assign _zz__zz__3_19_inner_macOut = ($signed(io_mulInput) * $signed(_3_19_inner_activation));
  assign _zz__zz__3_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_19_inner_macOut)) ? 16'h007f : _zz__3_19_inner_macOut_2);
  assign _zz__3_19_inner_macOut_2 = (($signed(_zz__3_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_19_inner_activation;
    end else begin
      io_macOut = _3_19_inner_macOut;
    end
  end

  assign _zz__3_19_inner_macOut = ($signed(_zz__zz__3_19_inner_macOut) + $signed(_zz__zz__3_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_19_inner_activation <= 8'h00;
      _3_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_19_inner_activation <= io_addInput;
      end else begin
        _3_19_inner_macOut <= _zz__3_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_114 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_18_inner_macOut;
  wire       [15:0]   _zz__zz__3_18_inner_macOut_1;
  wire       [15:0]   _zz__3_18_inner_macOut_1;
  wire       [15:0]   _zz__3_18_inner_macOut_2;
  reg        [7:0]    _3_18_inner_activation;
  reg        [7:0]    _3_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_18_inner_macOut;

  assign _zz__zz__3_18_inner_macOut = ($signed(io_mulInput) * $signed(_3_18_inner_activation));
  assign _zz__zz__3_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_18_inner_macOut)) ? 16'h007f : _zz__3_18_inner_macOut_2);
  assign _zz__3_18_inner_macOut_2 = (($signed(_zz__3_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_18_inner_activation;
    end else begin
      io_macOut = _3_18_inner_macOut;
    end
  end

  assign _zz__3_18_inner_macOut = ($signed(_zz__zz__3_18_inner_macOut) + $signed(_zz__zz__3_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_18_inner_activation <= 8'h00;
      _3_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_18_inner_activation <= io_addInput;
      end else begin
        _3_18_inner_macOut <= _zz__3_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_113 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_17_inner_macOut;
  wire       [15:0]   _zz__zz__3_17_inner_macOut_1;
  wire       [15:0]   _zz__3_17_inner_macOut_1;
  wire       [15:0]   _zz__3_17_inner_macOut_2;
  reg        [7:0]    _3_17_inner_activation;
  reg        [7:0]    _3_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_17_inner_macOut;

  assign _zz__zz__3_17_inner_macOut = ($signed(io_mulInput) * $signed(_3_17_inner_activation));
  assign _zz__zz__3_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_17_inner_macOut)) ? 16'h007f : _zz__3_17_inner_macOut_2);
  assign _zz__3_17_inner_macOut_2 = (($signed(_zz__3_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_17_inner_activation;
    end else begin
      io_macOut = _3_17_inner_macOut;
    end
  end

  assign _zz__3_17_inner_macOut = ($signed(_zz__zz__3_17_inner_macOut) + $signed(_zz__zz__3_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_17_inner_activation <= 8'h00;
      _3_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_17_inner_activation <= io_addInput;
      end else begin
        _3_17_inner_macOut <= _zz__3_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_112 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_16_inner_macOut;
  wire       [15:0]   _zz__zz__3_16_inner_macOut_1;
  wire       [15:0]   _zz__3_16_inner_macOut_1;
  wire       [15:0]   _zz__3_16_inner_macOut_2;
  reg        [7:0]    _3_16_inner_activation;
  reg        [7:0]    _3_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_16_inner_macOut;

  assign _zz__zz__3_16_inner_macOut = ($signed(io_mulInput) * $signed(_3_16_inner_activation));
  assign _zz__zz__3_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_16_inner_macOut)) ? 16'h007f : _zz__3_16_inner_macOut_2);
  assign _zz__3_16_inner_macOut_2 = (($signed(_zz__3_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_16_inner_activation;
    end else begin
      io_macOut = _3_16_inner_macOut;
    end
  end

  assign _zz__3_16_inner_macOut = ($signed(_zz__zz__3_16_inner_macOut) + $signed(_zz__zz__3_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_16_inner_activation <= 8'h00;
      _3_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_16_inner_activation <= io_addInput;
      end else begin
        _3_16_inner_macOut <= _zz__3_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_111 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_15_inner_macOut;
  wire       [15:0]   _zz__zz__3_15_inner_macOut_1;
  wire       [15:0]   _zz__3_15_inner_macOut_1;
  wire       [15:0]   _zz__3_15_inner_macOut_2;
  reg        [7:0]    _3_15_inner_activation;
  reg        [7:0]    _3_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_15_inner_macOut;

  assign _zz__zz__3_15_inner_macOut = ($signed(io_mulInput) * $signed(_3_15_inner_activation));
  assign _zz__zz__3_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_15_inner_macOut)) ? 16'h007f : _zz__3_15_inner_macOut_2);
  assign _zz__3_15_inner_macOut_2 = (($signed(_zz__3_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_15_inner_activation;
    end else begin
      io_macOut = _3_15_inner_macOut;
    end
  end

  assign _zz__3_15_inner_macOut = ($signed(_zz__zz__3_15_inner_macOut) + $signed(_zz__zz__3_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_15_inner_activation <= 8'h00;
      _3_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_15_inner_activation <= io_addInput;
      end else begin
        _3_15_inner_macOut <= _zz__3_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_110 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_14_inner_macOut;
  wire       [15:0]   _zz__zz__3_14_inner_macOut_1;
  wire       [15:0]   _zz__3_14_inner_macOut_1;
  wire       [15:0]   _zz__3_14_inner_macOut_2;
  reg        [7:0]    _3_14_inner_activation;
  reg        [7:0]    _3_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_14_inner_macOut;

  assign _zz__zz__3_14_inner_macOut = ($signed(io_mulInput) * $signed(_3_14_inner_activation));
  assign _zz__zz__3_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_14_inner_macOut)) ? 16'h007f : _zz__3_14_inner_macOut_2);
  assign _zz__3_14_inner_macOut_2 = (($signed(_zz__3_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_14_inner_activation;
    end else begin
      io_macOut = _3_14_inner_macOut;
    end
  end

  assign _zz__3_14_inner_macOut = ($signed(_zz__zz__3_14_inner_macOut) + $signed(_zz__zz__3_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_14_inner_activation <= 8'h00;
      _3_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_14_inner_activation <= io_addInput;
      end else begin
        _3_14_inner_macOut <= _zz__3_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_109 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_13_inner_macOut;
  wire       [15:0]   _zz__zz__3_13_inner_macOut_1;
  wire       [15:0]   _zz__3_13_inner_macOut_1;
  wire       [15:0]   _zz__3_13_inner_macOut_2;
  reg        [7:0]    _3_13_inner_activation;
  reg        [7:0]    _3_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_13_inner_macOut;

  assign _zz__zz__3_13_inner_macOut = ($signed(io_mulInput) * $signed(_3_13_inner_activation));
  assign _zz__zz__3_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_13_inner_macOut)) ? 16'h007f : _zz__3_13_inner_macOut_2);
  assign _zz__3_13_inner_macOut_2 = (($signed(_zz__3_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_13_inner_activation;
    end else begin
      io_macOut = _3_13_inner_macOut;
    end
  end

  assign _zz__3_13_inner_macOut = ($signed(_zz__zz__3_13_inner_macOut) + $signed(_zz__zz__3_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_13_inner_activation <= 8'h00;
      _3_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_13_inner_activation <= io_addInput;
      end else begin
        _3_13_inner_macOut <= _zz__3_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_108 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_12_inner_macOut;
  wire       [15:0]   _zz__zz__3_12_inner_macOut_1;
  wire       [15:0]   _zz__3_12_inner_macOut_1;
  wire       [15:0]   _zz__3_12_inner_macOut_2;
  reg        [7:0]    _3_12_inner_activation;
  reg        [7:0]    _3_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_12_inner_macOut;

  assign _zz__zz__3_12_inner_macOut = ($signed(io_mulInput) * $signed(_3_12_inner_activation));
  assign _zz__zz__3_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_12_inner_macOut)) ? 16'h007f : _zz__3_12_inner_macOut_2);
  assign _zz__3_12_inner_macOut_2 = (($signed(_zz__3_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_12_inner_activation;
    end else begin
      io_macOut = _3_12_inner_macOut;
    end
  end

  assign _zz__3_12_inner_macOut = ($signed(_zz__zz__3_12_inner_macOut) + $signed(_zz__zz__3_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_12_inner_activation <= 8'h00;
      _3_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_12_inner_activation <= io_addInput;
      end else begin
        _3_12_inner_macOut <= _zz__3_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_107 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_11_inner_macOut;
  wire       [15:0]   _zz__zz__3_11_inner_macOut_1;
  wire       [15:0]   _zz__3_11_inner_macOut_1;
  wire       [15:0]   _zz__3_11_inner_macOut_2;
  reg        [7:0]    _3_11_inner_activation;
  reg        [7:0]    _3_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_11_inner_macOut;

  assign _zz__zz__3_11_inner_macOut = ($signed(io_mulInput) * $signed(_3_11_inner_activation));
  assign _zz__zz__3_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_11_inner_macOut)) ? 16'h007f : _zz__3_11_inner_macOut_2);
  assign _zz__3_11_inner_macOut_2 = (($signed(_zz__3_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_11_inner_activation;
    end else begin
      io_macOut = _3_11_inner_macOut;
    end
  end

  assign _zz__3_11_inner_macOut = ($signed(_zz__zz__3_11_inner_macOut) + $signed(_zz__zz__3_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_11_inner_activation <= 8'h00;
      _3_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_11_inner_activation <= io_addInput;
      end else begin
        _3_11_inner_macOut <= _zz__3_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_106 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_10_inner_macOut;
  wire       [15:0]   _zz__zz__3_10_inner_macOut_1;
  wire       [15:0]   _zz__3_10_inner_macOut_1;
  wire       [15:0]   _zz__3_10_inner_macOut_2;
  reg        [7:0]    _3_10_inner_activation;
  reg        [7:0]    _3_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_10_inner_macOut;

  assign _zz__zz__3_10_inner_macOut = ($signed(io_mulInput) * $signed(_3_10_inner_activation));
  assign _zz__zz__3_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_10_inner_macOut)) ? 16'h007f : _zz__3_10_inner_macOut_2);
  assign _zz__3_10_inner_macOut_2 = (($signed(_zz__3_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_10_inner_activation;
    end else begin
      io_macOut = _3_10_inner_macOut;
    end
  end

  assign _zz__3_10_inner_macOut = ($signed(_zz__zz__3_10_inner_macOut) + $signed(_zz__zz__3_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_10_inner_activation <= 8'h00;
      _3_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_10_inner_activation <= io_addInput;
      end else begin
        _3_10_inner_macOut <= _zz__3_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_105 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_9_inner_macOut;
  wire       [15:0]   _zz__zz__3_9_inner_macOut_1;
  wire       [15:0]   _zz__3_9_inner_macOut_1;
  wire       [15:0]   _zz__3_9_inner_macOut_2;
  reg        [7:0]    _3_9_inner_activation;
  reg        [7:0]    _3_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_9_inner_macOut;

  assign _zz__zz__3_9_inner_macOut = ($signed(io_mulInput) * $signed(_3_9_inner_activation));
  assign _zz__zz__3_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_9_inner_macOut)) ? 16'h007f : _zz__3_9_inner_macOut_2);
  assign _zz__3_9_inner_macOut_2 = (($signed(_zz__3_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_9_inner_activation;
    end else begin
      io_macOut = _3_9_inner_macOut;
    end
  end

  assign _zz__3_9_inner_macOut = ($signed(_zz__zz__3_9_inner_macOut) + $signed(_zz__zz__3_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_9_inner_activation <= 8'h00;
      _3_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_9_inner_activation <= io_addInput;
      end else begin
        _3_9_inner_macOut <= _zz__3_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_104 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_8_inner_macOut;
  wire       [15:0]   _zz__zz__3_8_inner_macOut_1;
  wire       [15:0]   _zz__3_8_inner_macOut_1;
  wire       [15:0]   _zz__3_8_inner_macOut_2;
  reg        [7:0]    _3_8_inner_activation;
  reg        [7:0]    _3_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_8_inner_macOut;

  assign _zz__zz__3_8_inner_macOut = ($signed(io_mulInput) * $signed(_3_8_inner_activation));
  assign _zz__zz__3_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_8_inner_macOut)) ? 16'h007f : _zz__3_8_inner_macOut_2);
  assign _zz__3_8_inner_macOut_2 = (($signed(_zz__3_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_8_inner_activation;
    end else begin
      io_macOut = _3_8_inner_macOut;
    end
  end

  assign _zz__3_8_inner_macOut = ($signed(_zz__zz__3_8_inner_macOut) + $signed(_zz__zz__3_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_8_inner_activation <= 8'h00;
      _3_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_8_inner_activation <= io_addInput;
      end else begin
        _3_8_inner_macOut <= _zz__3_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_103 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_7_inner_macOut;
  wire       [15:0]   _zz__zz__3_7_inner_macOut_1;
  wire       [15:0]   _zz__3_7_inner_macOut_1;
  wire       [15:0]   _zz__3_7_inner_macOut_2;
  reg        [7:0]    _3_7_inner_activation;
  reg        [7:0]    _3_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_7_inner_macOut;

  assign _zz__zz__3_7_inner_macOut = ($signed(io_mulInput) * $signed(_3_7_inner_activation));
  assign _zz__zz__3_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_7_inner_macOut)) ? 16'h007f : _zz__3_7_inner_macOut_2);
  assign _zz__3_7_inner_macOut_2 = (($signed(_zz__3_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_7_inner_activation;
    end else begin
      io_macOut = _3_7_inner_macOut;
    end
  end

  assign _zz__3_7_inner_macOut = ($signed(_zz__zz__3_7_inner_macOut) + $signed(_zz__zz__3_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_7_inner_activation <= 8'h00;
      _3_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_7_inner_activation <= io_addInput;
      end else begin
        _3_7_inner_macOut <= _zz__3_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_102 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_6_inner_macOut;
  wire       [15:0]   _zz__zz__3_6_inner_macOut_1;
  wire       [15:0]   _zz__3_6_inner_macOut_1;
  wire       [15:0]   _zz__3_6_inner_macOut_2;
  reg        [7:0]    _3_6_inner_activation;
  reg        [7:0]    _3_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_6_inner_macOut;

  assign _zz__zz__3_6_inner_macOut = ($signed(io_mulInput) * $signed(_3_6_inner_activation));
  assign _zz__zz__3_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_6_inner_macOut)) ? 16'h007f : _zz__3_6_inner_macOut_2);
  assign _zz__3_6_inner_macOut_2 = (($signed(_zz__3_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_6_inner_activation;
    end else begin
      io_macOut = _3_6_inner_macOut;
    end
  end

  assign _zz__3_6_inner_macOut = ($signed(_zz__zz__3_6_inner_macOut) + $signed(_zz__zz__3_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_6_inner_activation <= 8'h00;
      _3_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_6_inner_activation <= io_addInput;
      end else begin
        _3_6_inner_macOut <= _zz__3_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_101 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_5_inner_macOut;
  wire       [15:0]   _zz__zz__3_5_inner_macOut_1;
  wire       [15:0]   _zz__3_5_inner_macOut_1;
  wire       [15:0]   _zz__3_5_inner_macOut_2;
  reg        [7:0]    _3_5_inner_activation;
  reg        [7:0]    _3_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_5_inner_macOut;

  assign _zz__zz__3_5_inner_macOut = ($signed(io_mulInput) * $signed(_3_5_inner_activation));
  assign _zz__zz__3_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_5_inner_macOut)) ? 16'h007f : _zz__3_5_inner_macOut_2);
  assign _zz__3_5_inner_macOut_2 = (($signed(_zz__3_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_5_inner_activation;
    end else begin
      io_macOut = _3_5_inner_macOut;
    end
  end

  assign _zz__3_5_inner_macOut = ($signed(_zz__zz__3_5_inner_macOut) + $signed(_zz__zz__3_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_5_inner_activation <= 8'h00;
      _3_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_5_inner_activation <= io_addInput;
      end else begin
        _3_5_inner_macOut <= _zz__3_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_100 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_4_inner_macOut;
  wire       [15:0]   _zz__zz__3_4_inner_macOut_1;
  wire       [15:0]   _zz__3_4_inner_macOut_1;
  wire       [15:0]   _zz__3_4_inner_macOut_2;
  reg        [7:0]    _3_4_inner_activation;
  reg        [7:0]    _3_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_4_inner_macOut;

  assign _zz__zz__3_4_inner_macOut = ($signed(io_mulInput) * $signed(_3_4_inner_activation));
  assign _zz__zz__3_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_4_inner_macOut)) ? 16'h007f : _zz__3_4_inner_macOut_2);
  assign _zz__3_4_inner_macOut_2 = (($signed(_zz__3_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_4_inner_activation;
    end else begin
      io_macOut = _3_4_inner_macOut;
    end
  end

  assign _zz__3_4_inner_macOut = ($signed(_zz__zz__3_4_inner_macOut) + $signed(_zz__zz__3_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_4_inner_activation <= 8'h00;
      _3_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_4_inner_activation <= io_addInput;
      end else begin
        _3_4_inner_macOut <= _zz__3_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_99 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_3_inner_macOut;
  wire       [15:0]   _zz__zz__3_3_inner_macOut_1;
  wire       [15:0]   _zz__3_3_inner_macOut_1;
  wire       [15:0]   _zz__3_3_inner_macOut_2;
  reg        [7:0]    _3_3_inner_activation;
  reg        [7:0]    _3_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_3_inner_macOut;

  assign _zz__zz__3_3_inner_macOut = ($signed(io_mulInput) * $signed(_3_3_inner_activation));
  assign _zz__zz__3_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_3_inner_macOut)) ? 16'h007f : _zz__3_3_inner_macOut_2);
  assign _zz__3_3_inner_macOut_2 = (($signed(_zz__3_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_3_inner_activation;
    end else begin
      io_macOut = _3_3_inner_macOut;
    end
  end

  assign _zz__3_3_inner_macOut = ($signed(_zz__zz__3_3_inner_macOut) + $signed(_zz__zz__3_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_3_inner_activation <= 8'h00;
      _3_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_3_inner_activation <= io_addInput;
      end else begin
        _3_3_inner_macOut <= _zz__3_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_98 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_2_inner_macOut;
  wire       [15:0]   _zz__zz__3_2_inner_macOut_1;
  wire       [15:0]   _zz__3_2_inner_macOut_1;
  wire       [15:0]   _zz__3_2_inner_macOut_2;
  reg        [7:0]    _3_2_inner_activation;
  reg        [7:0]    _3_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_2_inner_macOut;

  assign _zz__zz__3_2_inner_macOut = ($signed(io_mulInput) * $signed(_3_2_inner_activation));
  assign _zz__zz__3_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_2_inner_macOut)) ? 16'h007f : _zz__3_2_inner_macOut_2);
  assign _zz__3_2_inner_macOut_2 = (($signed(_zz__3_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_2_inner_activation;
    end else begin
      io_macOut = _3_2_inner_macOut;
    end
  end

  assign _zz__3_2_inner_macOut = ($signed(_zz__zz__3_2_inner_macOut) + $signed(_zz__zz__3_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_2_inner_activation <= 8'h00;
      _3_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_2_inner_activation <= io_addInput;
      end else begin
        _3_2_inner_macOut <= _zz__3_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_97 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_1_inner_macOut;
  wire       [15:0]   _zz__zz__3_1_inner_macOut_1;
  wire       [15:0]   _zz__3_1_inner_macOut_1;
  wire       [15:0]   _zz__3_1_inner_macOut_2;
  reg        [7:0]    _3_1_inner_activation;
  reg        [7:0]    _3_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_1_inner_macOut;

  assign _zz__zz__3_1_inner_macOut = ($signed(io_mulInput) * $signed(_3_1_inner_activation));
  assign _zz__zz__3_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_1_inner_macOut)) ? 16'h007f : _zz__3_1_inner_macOut_2);
  assign _zz__3_1_inner_macOut_2 = (($signed(_zz__3_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_1_inner_activation;
    end else begin
      io_macOut = _3_1_inner_macOut;
    end
  end

  assign _zz__3_1_inner_macOut = ($signed(_zz__zz__3_1_inner_macOut) + $signed(_zz__zz__3_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_1_inner_activation <= 8'h00;
      _3_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_1_inner_activation <= io_addInput;
      end else begin
        _3_1_inner_macOut <= _zz__3_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_96 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__3_0_inner_macOut;
  wire       [15:0]   _zz__zz__3_0_inner_macOut_1;
  wire       [15:0]   _zz__3_0_inner_macOut_1;
  wire       [15:0]   _zz__3_0_inner_macOut_2;
  reg        [7:0]    _3_0_inner_activation;
  reg        [7:0]    _3_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__3_0_inner_macOut;

  assign _zz__zz__3_0_inner_macOut = ($signed(io_mulInput) * $signed(_3_0_inner_activation));
  assign _zz__zz__3_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__3_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__3_0_inner_macOut)) ? 16'h007f : _zz__3_0_inner_macOut_2);
  assign _zz__3_0_inner_macOut_2 = (($signed(_zz__3_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__3_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _3_0_inner_activation;
    end else begin
      io_macOut = _3_0_inner_macOut;
    end
  end

  assign _zz__3_0_inner_macOut = ($signed(_zz__zz__3_0_inner_macOut) + $signed(_zz__zz__3_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _3_0_inner_activation <= 8'h00;
      _3_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _3_0_inner_activation <= io_addInput;
      end else begin
        _3_0_inner_macOut <= _zz__3_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_95 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_31_inner_macOut;
  wire       [15:0]   _zz__zz__2_31_inner_macOut_1;
  wire       [15:0]   _zz__2_31_inner_macOut_1;
  wire       [15:0]   _zz__2_31_inner_macOut_2;
  reg        [7:0]    _2_31_inner_activation;
  reg        [7:0]    _2_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_31_inner_macOut;

  assign _zz__zz__2_31_inner_macOut = ($signed(io_mulInput) * $signed(_2_31_inner_activation));
  assign _zz__zz__2_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_31_inner_macOut)) ? 16'h007f : _zz__2_31_inner_macOut_2);
  assign _zz__2_31_inner_macOut_2 = (($signed(_zz__2_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_31_inner_activation;
    end else begin
      io_macOut = _2_31_inner_macOut;
    end
  end

  assign _zz__2_31_inner_macOut = ($signed(_zz__zz__2_31_inner_macOut) + $signed(_zz__zz__2_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_31_inner_activation <= 8'h00;
      _2_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_31_inner_activation <= io_addInput;
      end else begin
        _2_31_inner_macOut <= _zz__2_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_94 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_30_inner_macOut;
  wire       [15:0]   _zz__zz__2_30_inner_macOut_1;
  wire       [15:0]   _zz__2_30_inner_macOut_1;
  wire       [15:0]   _zz__2_30_inner_macOut_2;
  reg        [7:0]    _2_30_inner_activation;
  reg        [7:0]    _2_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_30_inner_macOut;

  assign _zz__zz__2_30_inner_macOut = ($signed(io_mulInput) * $signed(_2_30_inner_activation));
  assign _zz__zz__2_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_30_inner_macOut)) ? 16'h007f : _zz__2_30_inner_macOut_2);
  assign _zz__2_30_inner_macOut_2 = (($signed(_zz__2_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_30_inner_activation;
    end else begin
      io_macOut = _2_30_inner_macOut;
    end
  end

  assign _zz__2_30_inner_macOut = ($signed(_zz__zz__2_30_inner_macOut) + $signed(_zz__zz__2_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_30_inner_activation <= 8'h00;
      _2_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_30_inner_activation <= io_addInput;
      end else begin
        _2_30_inner_macOut <= _zz__2_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_93 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_29_inner_macOut;
  wire       [15:0]   _zz__zz__2_29_inner_macOut_1;
  wire       [15:0]   _zz__2_29_inner_macOut_1;
  wire       [15:0]   _zz__2_29_inner_macOut_2;
  reg        [7:0]    _2_29_inner_activation;
  reg        [7:0]    _2_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_29_inner_macOut;

  assign _zz__zz__2_29_inner_macOut = ($signed(io_mulInput) * $signed(_2_29_inner_activation));
  assign _zz__zz__2_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_29_inner_macOut)) ? 16'h007f : _zz__2_29_inner_macOut_2);
  assign _zz__2_29_inner_macOut_2 = (($signed(_zz__2_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_29_inner_activation;
    end else begin
      io_macOut = _2_29_inner_macOut;
    end
  end

  assign _zz__2_29_inner_macOut = ($signed(_zz__zz__2_29_inner_macOut) + $signed(_zz__zz__2_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_29_inner_activation <= 8'h00;
      _2_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_29_inner_activation <= io_addInput;
      end else begin
        _2_29_inner_macOut <= _zz__2_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_92 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_28_inner_macOut;
  wire       [15:0]   _zz__zz__2_28_inner_macOut_1;
  wire       [15:0]   _zz__2_28_inner_macOut_1;
  wire       [15:0]   _zz__2_28_inner_macOut_2;
  reg        [7:0]    _2_28_inner_activation;
  reg        [7:0]    _2_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_28_inner_macOut;

  assign _zz__zz__2_28_inner_macOut = ($signed(io_mulInput) * $signed(_2_28_inner_activation));
  assign _zz__zz__2_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_28_inner_macOut)) ? 16'h007f : _zz__2_28_inner_macOut_2);
  assign _zz__2_28_inner_macOut_2 = (($signed(_zz__2_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_28_inner_activation;
    end else begin
      io_macOut = _2_28_inner_macOut;
    end
  end

  assign _zz__2_28_inner_macOut = ($signed(_zz__zz__2_28_inner_macOut) + $signed(_zz__zz__2_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_28_inner_activation <= 8'h00;
      _2_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_28_inner_activation <= io_addInput;
      end else begin
        _2_28_inner_macOut <= _zz__2_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_91 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_27_inner_macOut;
  wire       [15:0]   _zz__zz__2_27_inner_macOut_1;
  wire       [15:0]   _zz__2_27_inner_macOut_1;
  wire       [15:0]   _zz__2_27_inner_macOut_2;
  reg        [7:0]    _2_27_inner_activation;
  reg        [7:0]    _2_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_27_inner_macOut;

  assign _zz__zz__2_27_inner_macOut = ($signed(io_mulInput) * $signed(_2_27_inner_activation));
  assign _zz__zz__2_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_27_inner_macOut)) ? 16'h007f : _zz__2_27_inner_macOut_2);
  assign _zz__2_27_inner_macOut_2 = (($signed(_zz__2_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_27_inner_activation;
    end else begin
      io_macOut = _2_27_inner_macOut;
    end
  end

  assign _zz__2_27_inner_macOut = ($signed(_zz__zz__2_27_inner_macOut) + $signed(_zz__zz__2_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_27_inner_activation <= 8'h00;
      _2_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_27_inner_activation <= io_addInput;
      end else begin
        _2_27_inner_macOut <= _zz__2_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_90 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_26_inner_macOut;
  wire       [15:0]   _zz__zz__2_26_inner_macOut_1;
  wire       [15:0]   _zz__2_26_inner_macOut_1;
  wire       [15:0]   _zz__2_26_inner_macOut_2;
  reg        [7:0]    _2_26_inner_activation;
  reg        [7:0]    _2_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_26_inner_macOut;

  assign _zz__zz__2_26_inner_macOut = ($signed(io_mulInput) * $signed(_2_26_inner_activation));
  assign _zz__zz__2_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_26_inner_macOut)) ? 16'h007f : _zz__2_26_inner_macOut_2);
  assign _zz__2_26_inner_macOut_2 = (($signed(_zz__2_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_26_inner_activation;
    end else begin
      io_macOut = _2_26_inner_macOut;
    end
  end

  assign _zz__2_26_inner_macOut = ($signed(_zz__zz__2_26_inner_macOut) + $signed(_zz__zz__2_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_26_inner_activation <= 8'h00;
      _2_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_26_inner_activation <= io_addInput;
      end else begin
        _2_26_inner_macOut <= _zz__2_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_89 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_25_inner_macOut;
  wire       [15:0]   _zz__zz__2_25_inner_macOut_1;
  wire       [15:0]   _zz__2_25_inner_macOut_1;
  wire       [15:0]   _zz__2_25_inner_macOut_2;
  reg        [7:0]    _2_25_inner_activation;
  reg        [7:0]    _2_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_25_inner_macOut;

  assign _zz__zz__2_25_inner_macOut = ($signed(io_mulInput) * $signed(_2_25_inner_activation));
  assign _zz__zz__2_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_25_inner_macOut)) ? 16'h007f : _zz__2_25_inner_macOut_2);
  assign _zz__2_25_inner_macOut_2 = (($signed(_zz__2_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_25_inner_activation;
    end else begin
      io_macOut = _2_25_inner_macOut;
    end
  end

  assign _zz__2_25_inner_macOut = ($signed(_zz__zz__2_25_inner_macOut) + $signed(_zz__zz__2_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_25_inner_activation <= 8'h00;
      _2_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_25_inner_activation <= io_addInput;
      end else begin
        _2_25_inner_macOut <= _zz__2_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_88 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_24_inner_macOut;
  wire       [15:0]   _zz__zz__2_24_inner_macOut_1;
  wire       [15:0]   _zz__2_24_inner_macOut_1;
  wire       [15:0]   _zz__2_24_inner_macOut_2;
  reg        [7:0]    _2_24_inner_activation;
  reg        [7:0]    _2_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_24_inner_macOut;

  assign _zz__zz__2_24_inner_macOut = ($signed(io_mulInput) * $signed(_2_24_inner_activation));
  assign _zz__zz__2_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_24_inner_macOut)) ? 16'h007f : _zz__2_24_inner_macOut_2);
  assign _zz__2_24_inner_macOut_2 = (($signed(_zz__2_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_24_inner_activation;
    end else begin
      io_macOut = _2_24_inner_macOut;
    end
  end

  assign _zz__2_24_inner_macOut = ($signed(_zz__zz__2_24_inner_macOut) + $signed(_zz__zz__2_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_24_inner_activation <= 8'h00;
      _2_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_24_inner_activation <= io_addInput;
      end else begin
        _2_24_inner_macOut <= _zz__2_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_87 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_23_inner_macOut;
  wire       [15:0]   _zz__zz__2_23_inner_macOut_1;
  wire       [15:0]   _zz__2_23_inner_macOut_1;
  wire       [15:0]   _zz__2_23_inner_macOut_2;
  reg        [7:0]    _2_23_inner_activation;
  reg        [7:0]    _2_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_23_inner_macOut;

  assign _zz__zz__2_23_inner_macOut = ($signed(io_mulInput) * $signed(_2_23_inner_activation));
  assign _zz__zz__2_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_23_inner_macOut)) ? 16'h007f : _zz__2_23_inner_macOut_2);
  assign _zz__2_23_inner_macOut_2 = (($signed(_zz__2_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_23_inner_activation;
    end else begin
      io_macOut = _2_23_inner_macOut;
    end
  end

  assign _zz__2_23_inner_macOut = ($signed(_zz__zz__2_23_inner_macOut) + $signed(_zz__zz__2_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_23_inner_activation <= 8'h00;
      _2_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_23_inner_activation <= io_addInput;
      end else begin
        _2_23_inner_macOut <= _zz__2_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_86 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_22_inner_macOut;
  wire       [15:0]   _zz__zz__2_22_inner_macOut_1;
  wire       [15:0]   _zz__2_22_inner_macOut_1;
  wire       [15:0]   _zz__2_22_inner_macOut_2;
  reg        [7:0]    _2_22_inner_activation;
  reg        [7:0]    _2_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_22_inner_macOut;

  assign _zz__zz__2_22_inner_macOut = ($signed(io_mulInput) * $signed(_2_22_inner_activation));
  assign _zz__zz__2_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_22_inner_macOut)) ? 16'h007f : _zz__2_22_inner_macOut_2);
  assign _zz__2_22_inner_macOut_2 = (($signed(_zz__2_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_22_inner_activation;
    end else begin
      io_macOut = _2_22_inner_macOut;
    end
  end

  assign _zz__2_22_inner_macOut = ($signed(_zz__zz__2_22_inner_macOut) + $signed(_zz__zz__2_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_22_inner_activation <= 8'h00;
      _2_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_22_inner_activation <= io_addInput;
      end else begin
        _2_22_inner_macOut <= _zz__2_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_85 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_21_inner_macOut;
  wire       [15:0]   _zz__zz__2_21_inner_macOut_1;
  wire       [15:0]   _zz__2_21_inner_macOut_1;
  wire       [15:0]   _zz__2_21_inner_macOut_2;
  reg        [7:0]    _2_21_inner_activation;
  reg        [7:0]    _2_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_21_inner_macOut;

  assign _zz__zz__2_21_inner_macOut = ($signed(io_mulInput) * $signed(_2_21_inner_activation));
  assign _zz__zz__2_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_21_inner_macOut)) ? 16'h007f : _zz__2_21_inner_macOut_2);
  assign _zz__2_21_inner_macOut_2 = (($signed(_zz__2_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_21_inner_activation;
    end else begin
      io_macOut = _2_21_inner_macOut;
    end
  end

  assign _zz__2_21_inner_macOut = ($signed(_zz__zz__2_21_inner_macOut) + $signed(_zz__zz__2_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_21_inner_activation <= 8'h00;
      _2_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_21_inner_activation <= io_addInput;
      end else begin
        _2_21_inner_macOut <= _zz__2_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_84 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_20_inner_macOut;
  wire       [15:0]   _zz__zz__2_20_inner_macOut_1;
  wire       [15:0]   _zz__2_20_inner_macOut_1;
  wire       [15:0]   _zz__2_20_inner_macOut_2;
  reg        [7:0]    _2_20_inner_activation;
  reg        [7:0]    _2_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_20_inner_macOut;

  assign _zz__zz__2_20_inner_macOut = ($signed(io_mulInput) * $signed(_2_20_inner_activation));
  assign _zz__zz__2_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_20_inner_macOut)) ? 16'h007f : _zz__2_20_inner_macOut_2);
  assign _zz__2_20_inner_macOut_2 = (($signed(_zz__2_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_20_inner_activation;
    end else begin
      io_macOut = _2_20_inner_macOut;
    end
  end

  assign _zz__2_20_inner_macOut = ($signed(_zz__zz__2_20_inner_macOut) + $signed(_zz__zz__2_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_20_inner_activation <= 8'h00;
      _2_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_20_inner_activation <= io_addInput;
      end else begin
        _2_20_inner_macOut <= _zz__2_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_83 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_19_inner_macOut;
  wire       [15:0]   _zz__zz__2_19_inner_macOut_1;
  wire       [15:0]   _zz__2_19_inner_macOut_1;
  wire       [15:0]   _zz__2_19_inner_macOut_2;
  reg        [7:0]    _2_19_inner_activation;
  reg        [7:0]    _2_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_19_inner_macOut;

  assign _zz__zz__2_19_inner_macOut = ($signed(io_mulInput) * $signed(_2_19_inner_activation));
  assign _zz__zz__2_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_19_inner_macOut)) ? 16'h007f : _zz__2_19_inner_macOut_2);
  assign _zz__2_19_inner_macOut_2 = (($signed(_zz__2_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_19_inner_activation;
    end else begin
      io_macOut = _2_19_inner_macOut;
    end
  end

  assign _zz__2_19_inner_macOut = ($signed(_zz__zz__2_19_inner_macOut) + $signed(_zz__zz__2_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_19_inner_activation <= 8'h00;
      _2_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_19_inner_activation <= io_addInput;
      end else begin
        _2_19_inner_macOut <= _zz__2_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_82 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_18_inner_macOut;
  wire       [15:0]   _zz__zz__2_18_inner_macOut_1;
  wire       [15:0]   _zz__2_18_inner_macOut_1;
  wire       [15:0]   _zz__2_18_inner_macOut_2;
  reg        [7:0]    _2_18_inner_activation;
  reg        [7:0]    _2_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_18_inner_macOut;

  assign _zz__zz__2_18_inner_macOut = ($signed(io_mulInput) * $signed(_2_18_inner_activation));
  assign _zz__zz__2_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_18_inner_macOut)) ? 16'h007f : _zz__2_18_inner_macOut_2);
  assign _zz__2_18_inner_macOut_2 = (($signed(_zz__2_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_18_inner_activation;
    end else begin
      io_macOut = _2_18_inner_macOut;
    end
  end

  assign _zz__2_18_inner_macOut = ($signed(_zz__zz__2_18_inner_macOut) + $signed(_zz__zz__2_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_18_inner_activation <= 8'h00;
      _2_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_18_inner_activation <= io_addInput;
      end else begin
        _2_18_inner_macOut <= _zz__2_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_81 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_17_inner_macOut;
  wire       [15:0]   _zz__zz__2_17_inner_macOut_1;
  wire       [15:0]   _zz__2_17_inner_macOut_1;
  wire       [15:0]   _zz__2_17_inner_macOut_2;
  reg        [7:0]    _2_17_inner_activation;
  reg        [7:0]    _2_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_17_inner_macOut;

  assign _zz__zz__2_17_inner_macOut = ($signed(io_mulInput) * $signed(_2_17_inner_activation));
  assign _zz__zz__2_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_17_inner_macOut)) ? 16'h007f : _zz__2_17_inner_macOut_2);
  assign _zz__2_17_inner_macOut_2 = (($signed(_zz__2_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_17_inner_activation;
    end else begin
      io_macOut = _2_17_inner_macOut;
    end
  end

  assign _zz__2_17_inner_macOut = ($signed(_zz__zz__2_17_inner_macOut) + $signed(_zz__zz__2_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_17_inner_activation <= 8'h00;
      _2_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_17_inner_activation <= io_addInput;
      end else begin
        _2_17_inner_macOut <= _zz__2_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_80 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_16_inner_macOut;
  wire       [15:0]   _zz__zz__2_16_inner_macOut_1;
  wire       [15:0]   _zz__2_16_inner_macOut_1;
  wire       [15:0]   _zz__2_16_inner_macOut_2;
  reg        [7:0]    _2_16_inner_activation;
  reg        [7:0]    _2_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_16_inner_macOut;

  assign _zz__zz__2_16_inner_macOut = ($signed(io_mulInput) * $signed(_2_16_inner_activation));
  assign _zz__zz__2_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_16_inner_macOut)) ? 16'h007f : _zz__2_16_inner_macOut_2);
  assign _zz__2_16_inner_macOut_2 = (($signed(_zz__2_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_16_inner_activation;
    end else begin
      io_macOut = _2_16_inner_macOut;
    end
  end

  assign _zz__2_16_inner_macOut = ($signed(_zz__zz__2_16_inner_macOut) + $signed(_zz__zz__2_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_16_inner_activation <= 8'h00;
      _2_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_16_inner_activation <= io_addInput;
      end else begin
        _2_16_inner_macOut <= _zz__2_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_79 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_15_inner_macOut;
  wire       [15:0]   _zz__zz__2_15_inner_macOut_1;
  wire       [15:0]   _zz__2_15_inner_macOut_1;
  wire       [15:0]   _zz__2_15_inner_macOut_2;
  reg        [7:0]    _2_15_inner_activation;
  reg        [7:0]    _2_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_15_inner_macOut;

  assign _zz__zz__2_15_inner_macOut = ($signed(io_mulInput) * $signed(_2_15_inner_activation));
  assign _zz__zz__2_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_15_inner_macOut)) ? 16'h007f : _zz__2_15_inner_macOut_2);
  assign _zz__2_15_inner_macOut_2 = (($signed(_zz__2_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_15_inner_activation;
    end else begin
      io_macOut = _2_15_inner_macOut;
    end
  end

  assign _zz__2_15_inner_macOut = ($signed(_zz__zz__2_15_inner_macOut) + $signed(_zz__zz__2_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_15_inner_activation <= 8'h00;
      _2_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_15_inner_activation <= io_addInput;
      end else begin
        _2_15_inner_macOut <= _zz__2_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_78 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_14_inner_macOut;
  wire       [15:0]   _zz__zz__2_14_inner_macOut_1;
  wire       [15:0]   _zz__2_14_inner_macOut_1;
  wire       [15:0]   _zz__2_14_inner_macOut_2;
  reg        [7:0]    _2_14_inner_activation;
  reg        [7:0]    _2_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_14_inner_macOut;

  assign _zz__zz__2_14_inner_macOut = ($signed(io_mulInput) * $signed(_2_14_inner_activation));
  assign _zz__zz__2_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_14_inner_macOut)) ? 16'h007f : _zz__2_14_inner_macOut_2);
  assign _zz__2_14_inner_macOut_2 = (($signed(_zz__2_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_14_inner_activation;
    end else begin
      io_macOut = _2_14_inner_macOut;
    end
  end

  assign _zz__2_14_inner_macOut = ($signed(_zz__zz__2_14_inner_macOut) + $signed(_zz__zz__2_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_14_inner_activation <= 8'h00;
      _2_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_14_inner_activation <= io_addInput;
      end else begin
        _2_14_inner_macOut <= _zz__2_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_77 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_13_inner_macOut;
  wire       [15:0]   _zz__zz__2_13_inner_macOut_1;
  wire       [15:0]   _zz__2_13_inner_macOut_1;
  wire       [15:0]   _zz__2_13_inner_macOut_2;
  reg        [7:0]    _2_13_inner_activation;
  reg        [7:0]    _2_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_13_inner_macOut;

  assign _zz__zz__2_13_inner_macOut = ($signed(io_mulInput) * $signed(_2_13_inner_activation));
  assign _zz__zz__2_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_13_inner_macOut)) ? 16'h007f : _zz__2_13_inner_macOut_2);
  assign _zz__2_13_inner_macOut_2 = (($signed(_zz__2_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_13_inner_activation;
    end else begin
      io_macOut = _2_13_inner_macOut;
    end
  end

  assign _zz__2_13_inner_macOut = ($signed(_zz__zz__2_13_inner_macOut) + $signed(_zz__zz__2_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_13_inner_activation <= 8'h00;
      _2_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_13_inner_activation <= io_addInput;
      end else begin
        _2_13_inner_macOut <= _zz__2_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_76 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_12_inner_macOut;
  wire       [15:0]   _zz__zz__2_12_inner_macOut_1;
  wire       [15:0]   _zz__2_12_inner_macOut_1;
  wire       [15:0]   _zz__2_12_inner_macOut_2;
  reg        [7:0]    _2_12_inner_activation;
  reg        [7:0]    _2_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_12_inner_macOut;

  assign _zz__zz__2_12_inner_macOut = ($signed(io_mulInput) * $signed(_2_12_inner_activation));
  assign _zz__zz__2_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_12_inner_macOut)) ? 16'h007f : _zz__2_12_inner_macOut_2);
  assign _zz__2_12_inner_macOut_2 = (($signed(_zz__2_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_12_inner_activation;
    end else begin
      io_macOut = _2_12_inner_macOut;
    end
  end

  assign _zz__2_12_inner_macOut = ($signed(_zz__zz__2_12_inner_macOut) + $signed(_zz__zz__2_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_12_inner_activation <= 8'h00;
      _2_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_12_inner_activation <= io_addInput;
      end else begin
        _2_12_inner_macOut <= _zz__2_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_75 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_11_inner_macOut;
  wire       [15:0]   _zz__zz__2_11_inner_macOut_1;
  wire       [15:0]   _zz__2_11_inner_macOut_1;
  wire       [15:0]   _zz__2_11_inner_macOut_2;
  reg        [7:0]    _2_11_inner_activation;
  reg        [7:0]    _2_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_11_inner_macOut;

  assign _zz__zz__2_11_inner_macOut = ($signed(io_mulInput) * $signed(_2_11_inner_activation));
  assign _zz__zz__2_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_11_inner_macOut)) ? 16'h007f : _zz__2_11_inner_macOut_2);
  assign _zz__2_11_inner_macOut_2 = (($signed(_zz__2_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_11_inner_activation;
    end else begin
      io_macOut = _2_11_inner_macOut;
    end
  end

  assign _zz__2_11_inner_macOut = ($signed(_zz__zz__2_11_inner_macOut) + $signed(_zz__zz__2_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_11_inner_activation <= 8'h00;
      _2_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_11_inner_activation <= io_addInput;
      end else begin
        _2_11_inner_macOut <= _zz__2_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_74 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_10_inner_macOut;
  wire       [15:0]   _zz__zz__2_10_inner_macOut_1;
  wire       [15:0]   _zz__2_10_inner_macOut_1;
  wire       [15:0]   _zz__2_10_inner_macOut_2;
  reg        [7:0]    _2_10_inner_activation;
  reg        [7:0]    _2_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_10_inner_macOut;

  assign _zz__zz__2_10_inner_macOut = ($signed(io_mulInput) * $signed(_2_10_inner_activation));
  assign _zz__zz__2_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_10_inner_macOut)) ? 16'h007f : _zz__2_10_inner_macOut_2);
  assign _zz__2_10_inner_macOut_2 = (($signed(_zz__2_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_10_inner_activation;
    end else begin
      io_macOut = _2_10_inner_macOut;
    end
  end

  assign _zz__2_10_inner_macOut = ($signed(_zz__zz__2_10_inner_macOut) + $signed(_zz__zz__2_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_10_inner_activation <= 8'h00;
      _2_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_10_inner_activation <= io_addInput;
      end else begin
        _2_10_inner_macOut <= _zz__2_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_73 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_9_inner_macOut;
  wire       [15:0]   _zz__zz__2_9_inner_macOut_1;
  wire       [15:0]   _zz__2_9_inner_macOut_1;
  wire       [15:0]   _zz__2_9_inner_macOut_2;
  reg        [7:0]    _2_9_inner_activation;
  reg        [7:0]    _2_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_9_inner_macOut;

  assign _zz__zz__2_9_inner_macOut = ($signed(io_mulInput) * $signed(_2_9_inner_activation));
  assign _zz__zz__2_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_9_inner_macOut)) ? 16'h007f : _zz__2_9_inner_macOut_2);
  assign _zz__2_9_inner_macOut_2 = (($signed(_zz__2_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_9_inner_activation;
    end else begin
      io_macOut = _2_9_inner_macOut;
    end
  end

  assign _zz__2_9_inner_macOut = ($signed(_zz__zz__2_9_inner_macOut) + $signed(_zz__zz__2_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_9_inner_activation <= 8'h00;
      _2_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_9_inner_activation <= io_addInput;
      end else begin
        _2_9_inner_macOut <= _zz__2_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_72 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_8_inner_macOut;
  wire       [15:0]   _zz__zz__2_8_inner_macOut_1;
  wire       [15:0]   _zz__2_8_inner_macOut_1;
  wire       [15:0]   _zz__2_8_inner_macOut_2;
  reg        [7:0]    _2_8_inner_activation;
  reg        [7:0]    _2_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_8_inner_macOut;

  assign _zz__zz__2_8_inner_macOut = ($signed(io_mulInput) * $signed(_2_8_inner_activation));
  assign _zz__zz__2_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_8_inner_macOut)) ? 16'h007f : _zz__2_8_inner_macOut_2);
  assign _zz__2_8_inner_macOut_2 = (($signed(_zz__2_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_8_inner_activation;
    end else begin
      io_macOut = _2_8_inner_macOut;
    end
  end

  assign _zz__2_8_inner_macOut = ($signed(_zz__zz__2_8_inner_macOut) + $signed(_zz__zz__2_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_8_inner_activation <= 8'h00;
      _2_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_8_inner_activation <= io_addInput;
      end else begin
        _2_8_inner_macOut <= _zz__2_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_71 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_7_inner_macOut;
  wire       [15:0]   _zz__zz__2_7_inner_macOut_1;
  wire       [15:0]   _zz__2_7_inner_macOut_1;
  wire       [15:0]   _zz__2_7_inner_macOut_2;
  reg        [7:0]    _2_7_inner_activation;
  reg        [7:0]    _2_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_7_inner_macOut;

  assign _zz__zz__2_7_inner_macOut = ($signed(io_mulInput) * $signed(_2_7_inner_activation));
  assign _zz__zz__2_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_7_inner_macOut)) ? 16'h007f : _zz__2_7_inner_macOut_2);
  assign _zz__2_7_inner_macOut_2 = (($signed(_zz__2_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_7_inner_activation;
    end else begin
      io_macOut = _2_7_inner_macOut;
    end
  end

  assign _zz__2_7_inner_macOut = ($signed(_zz__zz__2_7_inner_macOut) + $signed(_zz__zz__2_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_7_inner_activation <= 8'h00;
      _2_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_7_inner_activation <= io_addInput;
      end else begin
        _2_7_inner_macOut <= _zz__2_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_70 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_6_inner_macOut;
  wire       [15:0]   _zz__zz__2_6_inner_macOut_1;
  wire       [15:0]   _zz__2_6_inner_macOut_1;
  wire       [15:0]   _zz__2_6_inner_macOut_2;
  reg        [7:0]    _2_6_inner_activation;
  reg        [7:0]    _2_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_6_inner_macOut;

  assign _zz__zz__2_6_inner_macOut = ($signed(io_mulInput) * $signed(_2_6_inner_activation));
  assign _zz__zz__2_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_6_inner_macOut)) ? 16'h007f : _zz__2_6_inner_macOut_2);
  assign _zz__2_6_inner_macOut_2 = (($signed(_zz__2_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_6_inner_activation;
    end else begin
      io_macOut = _2_6_inner_macOut;
    end
  end

  assign _zz__2_6_inner_macOut = ($signed(_zz__zz__2_6_inner_macOut) + $signed(_zz__zz__2_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_6_inner_activation <= 8'h00;
      _2_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_6_inner_activation <= io_addInput;
      end else begin
        _2_6_inner_macOut <= _zz__2_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_69 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_5_inner_macOut;
  wire       [15:0]   _zz__zz__2_5_inner_macOut_1;
  wire       [15:0]   _zz__2_5_inner_macOut_1;
  wire       [15:0]   _zz__2_5_inner_macOut_2;
  reg        [7:0]    _2_5_inner_activation;
  reg        [7:0]    _2_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_5_inner_macOut;

  assign _zz__zz__2_5_inner_macOut = ($signed(io_mulInput) * $signed(_2_5_inner_activation));
  assign _zz__zz__2_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_5_inner_macOut)) ? 16'h007f : _zz__2_5_inner_macOut_2);
  assign _zz__2_5_inner_macOut_2 = (($signed(_zz__2_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_5_inner_activation;
    end else begin
      io_macOut = _2_5_inner_macOut;
    end
  end

  assign _zz__2_5_inner_macOut = ($signed(_zz__zz__2_5_inner_macOut) + $signed(_zz__zz__2_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_5_inner_activation <= 8'h00;
      _2_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_5_inner_activation <= io_addInput;
      end else begin
        _2_5_inner_macOut <= _zz__2_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_68 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_4_inner_macOut;
  wire       [15:0]   _zz__zz__2_4_inner_macOut_1;
  wire       [15:0]   _zz__2_4_inner_macOut_1;
  wire       [15:0]   _zz__2_4_inner_macOut_2;
  reg        [7:0]    _2_4_inner_activation;
  reg        [7:0]    _2_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_4_inner_macOut;

  assign _zz__zz__2_4_inner_macOut = ($signed(io_mulInput) * $signed(_2_4_inner_activation));
  assign _zz__zz__2_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_4_inner_macOut)) ? 16'h007f : _zz__2_4_inner_macOut_2);
  assign _zz__2_4_inner_macOut_2 = (($signed(_zz__2_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_4_inner_activation;
    end else begin
      io_macOut = _2_4_inner_macOut;
    end
  end

  assign _zz__2_4_inner_macOut = ($signed(_zz__zz__2_4_inner_macOut) + $signed(_zz__zz__2_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_4_inner_activation <= 8'h00;
      _2_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_4_inner_activation <= io_addInput;
      end else begin
        _2_4_inner_macOut <= _zz__2_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_67 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_3_inner_macOut;
  wire       [15:0]   _zz__zz__2_3_inner_macOut_1;
  wire       [15:0]   _zz__2_3_inner_macOut_1;
  wire       [15:0]   _zz__2_3_inner_macOut_2;
  reg        [7:0]    _2_3_inner_activation;
  reg        [7:0]    _2_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_3_inner_macOut;

  assign _zz__zz__2_3_inner_macOut = ($signed(io_mulInput) * $signed(_2_3_inner_activation));
  assign _zz__zz__2_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_3_inner_macOut)) ? 16'h007f : _zz__2_3_inner_macOut_2);
  assign _zz__2_3_inner_macOut_2 = (($signed(_zz__2_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_3_inner_activation;
    end else begin
      io_macOut = _2_3_inner_macOut;
    end
  end

  assign _zz__2_3_inner_macOut = ($signed(_zz__zz__2_3_inner_macOut) + $signed(_zz__zz__2_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_3_inner_activation <= 8'h00;
      _2_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_3_inner_activation <= io_addInput;
      end else begin
        _2_3_inner_macOut <= _zz__2_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_66 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_2_inner_macOut;
  wire       [15:0]   _zz__zz__2_2_inner_macOut_1;
  wire       [15:0]   _zz__2_2_inner_macOut_1;
  wire       [15:0]   _zz__2_2_inner_macOut_2;
  reg        [7:0]    _2_2_inner_activation;
  reg        [7:0]    _2_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_2_inner_macOut;

  assign _zz__zz__2_2_inner_macOut = ($signed(io_mulInput) * $signed(_2_2_inner_activation));
  assign _zz__zz__2_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_2_inner_macOut)) ? 16'h007f : _zz__2_2_inner_macOut_2);
  assign _zz__2_2_inner_macOut_2 = (($signed(_zz__2_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_2_inner_activation;
    end else begin
      io_macOut = _2_2_inner_macOut;
    end
  end

  assign _zz__2_2_inner_macOut = ($signed(_zz__zz__2_2_inner_macOut) + $signed(_zz__zz__2_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_2_inner_activation <= 8'h00;
      _2_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_2_inner_activation <= io_addInput;
      end else begin
        _2_2_inner_macOut <= _zz__2_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_65 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_1_inner_macOut;
  wire       [15:0]   _zz__zz__2_1_inner_macOut_1;
  wire       [15:0]   _zz__2_1_inner_macOut_1;
  wire       [15:0]   _zz__2_1_inner_macOut_2;
  reg        [7:0]    _2_1_inner_activation;
  reg        [7:0]    _2_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_1_inner_macOut;

  assign _zz__zz__2_1_inner_macOut = ($signed(io_mulInput) * $signed(_2_1_inner_activation));
  assign _zz__zz__2_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_1_inner_macOut)) ? 16'h007f : _zz__2_1_inner_macOut_2);
  assign _zz__2_1_inner_macOut_2 = (($signed(_zz__2_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_1_inner_activation;
    end else begin
      io_macOut = _2_1_inner_macOut;
    end
  end

  assign _zz__2_1_inner_macOut = ($signed(_zz__zz__2_1_inner_macOut) + $signed(_zz__zz__2_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_1_inner_activation <= 8'h00;
      _2_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_1_inner_activation <= io_addInput;
      end else begin
        _2_1_inner_macOut <= _zz__2_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_64 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__2_0_inner_macOut;
  wire       [15:0]   _zz__zz__2_0_inner_macOut_1;
  wire       [15:0]   _zz__2_0_inner_macOut_1;
  wire       [15:0]   _zz__2_0_inner_macOut_2;
  reg        [7:0]    _2_0_inner_activation;
  reg        [7:0]    _2_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__2_0_inner_macOut;

  assign _zz__zz__2_0_inner_macOut = ($signed(io_mulInput) * $signed(_2_0_inner_activation));
  assign _zz__zz__2_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__2_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__2_0_inner_macOut)) ? 16'h007f : _zz__2_0_inner_macOut_2);
  assign _zz__2_0_inner_macOut_2 = (($signed(_zz__2_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__2_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _2_0_inner_activation;
    end else begin
      io_macOut = _2_0_inner_macOut;
    end
  end

  assign _zz__2_0_inner_macOut = ($signed(_zz__zz__2_0_inner_macOut) + $signed(_zz__zz__2_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _2_0_inner_activation <= 8'h00;
      _2_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _2_0_inner_activation <= io_addInput;
      end else begin
        _2_0_inner_macOut <= _zz__2_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_63 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_31_inner_macOut;
  wire       [15:0]   _zz__zz__1_31_inner_macOut_1;
  wire       [15:0]   _zz__1_31_inner_macOut_1;
  wire       [15:0]   _zz__1_31_inner_macOut_2;
  reg        [7:0]    _1_31_inner_activation;
  reg        [7:0]    _1_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_31_inner_macOut;

  assign _zz__zz__1_31_inner_macOut = ($signed(io_mulInput) * $signed(_1_31_inner_activation));
  assign _zz__zz__1_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_31_inner_macOut)) ? 16'h007f : _zz__1_31_inner_macOut_2);
  assign _zz__1_31_inner_macOut_2 = (($signed(_zz__1_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_31_inner_activation;
    end else begin
      io_macOut = _1_31_inner_macOut;
    end
  end

  assign _zz__1_31_inner_macOut = ($signed(_zz__zz__1_31_inner_macOut) + $signed(_zz__zz__1_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_31_inner_activation <= 8'h00;
      _1_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_31_inner_activation <= io_addInput;
      end else begin
        _1_31_inner_macOut <= _zz__1_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_62 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_30_inner_macOut;
  wire       [15:0]   _zz__zz__1_30_inner_macOut_1;
  wire       [15:0]   _zz__1_30_inner_macOut_1;
  wire       [15:0]   _zz__1_30_inner_macOut_2;
  reg        [7:0]    _1_30_inner_activation;
  reg        [7:0]    _1_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_30_inner_macOut;

  assign _zz__zz__1_30_inner_macOut = ($signed(io_mulInput) * $signed(_1_30_inner_activation));
  assign _zz__zz__1_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_30_inner_macOut)) ? 16'h007f : _zz__1_30_inner_macOut_2);
  assign _zz__1_30_inner_macOut_2 = (($signed(_zz__1_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_30_inner_activation;
    end else begin
      io_macOut = _1_30_inner_macOut;
    end
  end

  assign _zz__1_30_inner_macOut = ($signed(_zz__zz__1_30_inner_macOut) + $signed(_zz__zz__1_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_30_inner_activation <= 8'h00;
      _1_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_30_inner_activation <= io_addInput;
      end else begin
        _1_30_inner_macOut <= _zz__1_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_61 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_29_inner_macOut;
  wire       [15:0]   _zz__zz__1_29_inner_macOut_1;
  wire       [15:0]   _zz__1_29_inner_macOut_1;
  wire       [15:0]   _zz__1_29_inner_macOut_2;
  reg        [7:0]    _1_29_inner_activation;
  reg        [7:0]    _1_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_29_inner_macOut;

  assign _zz__zz__1_29_inner_macOut = ($signed(io_mulInput) * $signed(_1_29_inner_activation));
  assign _zz__zz__1_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_29_inner_macOut)) ? 16'h007f : _zz__1_29_inner_macOut_2);
  assign _zz__1_29_inner_macOut_2 = (($signed(_zz__1_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_29_inner_activation;
    end else begin
      io_macOut = _1_29_inner_macOut;
    end
  end

  assign _zz__1_29_inner_macOut = ($signed(_zz__zz__1_29_inner_macOut) + $signed(_zz__zz__1_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_29_inner_activation <= 8'h00;
      _1_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_29_inner_activation <= io_addInput;
      end else begin
        _1_29_inner_macOut <= _zz__1_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_60 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_28_inner_macOut;
  wire       [15:0]   _zz__zz__1_28_inner_macOut_1;
  wire       [15:0]   _zz__1_28_inner_macOut_1;
  wire       [15:0]   _zz__1_28_inner_macOut_2;
  reg        [7:0]    _1_28_inner_activation;
  reg        [7:0]    _1_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_28_inner_macOut;

  assign _zz__zz__1_28_inner_macOut = ($signed(io_mulInput) * $signed(_1_28_inner_activation));
  assign _zz__zz__1_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_28_inner_macOut)) ? 16'h007f : _zz__1_28_inner_macOut_2);
  assign _zz__1_28_inner_macOut_2 = (($signed(_zz__1_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_28_inner_activation;
    end else begin
      io_macOut = _1_28_inner_macOut;
    end
  end

  assign _zz__1_28_inner_macOut = ($signed(_zz__zz__1_28_inner_macOut) + $signed(_zz__zz__1_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_28_inner_activation <= 8'h00;
      _1_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_28_inner_activation <= io_addInput;
      end else begin
        _1_28_inner_macOut <= _zz__1_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_59 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_27_inner_macOut;
  wire       [15:0]   _zz__zz__1_27_inner_macOut_1;
  wire       [15:0]   _zz__1_27_inner_macOut_1;
  wire       [15:0]   _zz__1_27_inner_macOut_2;
  reg        [7:0]    _1_27_inner_activation;
  reg        [7:0]    _1_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_27_inner_macOut;

  assign _zz__zz__1_27_inner_macOut = ($signed(io_mulInput) * $signed(_1_27_inner_activation));
  assign _zz__zz__1_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_27_inner_macOut)) ? 16'h007f : _zz__1_27_inner_macOut_2);
  assign _zz__1_27_inner_macOut_2 = (($signed(_zz__1_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_27_inner_activation;
    end else begin
      io_macOut = _1_27_inner_macOut;
    end
  end

  assign _zz__1_27_inner_macOut = ($signed(_zz__zz__1_27_inner_macOut) + $signed(_zz__zz__1_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_27_inner_activation <= 8'h00;
      _1_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_27_inner_activation <= io_addInput;
      end else begin
        _1_27_inner_macOut <= _zz__1_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_58 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_26_inner_macOut;
  wire       [15:0]   _zz__zz__1_26_inner_macOut_1;
  wire       [15:0]   _zz__1_26_inner_macOut_1;
  wire       [15:0]   _zz__1_26_inner_macOut_2;
  reg        [7:0]    _1_26_inner_activation;
  reg        [7:0]    _1_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_26_inner_macOut;

  assign _zz__zz__1_26_inner_macOut = ($signed(io_mulInput) * $signed(_1_26_inner_activation));
  assign _zz__zz__1_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_26_inner_macOut)) ? 16'h007f : _zz__1_26_inner_macOut_2);
  assign _zz__1_26_inner_macOut_2 = (($signed(_zz__1_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_26_inner_activation;
    end else begin
      io_macOut = _1_26_inner_macOut;
    end
  end

  assign _zz__1_26_inner_macOut = ($signed(_zz__zz__1_26_inner_macOut) + $signed(_zz__zz__1_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_26_inner_activation <= 8'h00;
      _1_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_26_inner_activation <= io_addInput;
      end else begin
        _1_26_inner_macOut <= _zz__1_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_57 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_25_inner_macOut;
  wire       [15:0]   _zz__zz__1_25_inner_macOut_1;
  wire       [15:0]   _zz__1_25_inner_macOut_1;
  wire       [15:0]   _zz__1_25_inner_macOut_2;
  reg        [7:0]    _1_25_inner_activation;
  reg        [7:0]    _1_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_25_inner_macOut;

  assign _zz__zz__1_25_inner_macOut = ($signed(io_mulInput) * $signed(_1_25_inner_activation));
  assign _zz__zz__1_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_25_inner_macOut)) ? 16'h007f : _zz__1_25_inner_macOut_2);
  assign _zz__1_25_inner_macOut_2 = (($signed(_zz__1_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_25_inner_activation;
    end else begin
      io_macOut = _1_25_inner_macOut;
    end
  end

  assign _zz__1_25_inner_macOut = ($signed(_zz__zz__1_25_inner_macOut) + $signed(_zz__zz__1_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_25_inner_activation <= 8'h00;
      _1_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_25_inner_activation <= io_addInput;
      end else begin
        _1_25_inner_macOut <= _zz__1_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_56 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_24_inner_macOut;
  wire       [15:0]   _zz__zz__1_24_inner_macOut_1;
  wire       [15:0]   _zz__1_24_inner_macOut_1;
  wire       [15:0]   _zz__1_24_inner_macOut_2;
  reg        [7:0]    _1_24_inner_activation;
  reg        [7:0]    _1_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_24_inner_macOut;

  assign _zz__zz__1_24_inner_macOut = ($signed(io_mulInput) * $signed(_1_24_inner_activation));
  assign _zz__zz__1_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_24_inner_macOut)) ? 16'h007f : _zz__1_24_inner_macOut_2);
  assign _zz__1_24_inner_macOut_2 = (($signed(_zz__1_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_24_inner_activation;
    end else begin
      io_macOut = _1_24_inner_macOut;
    end
  end

  assign _zz__1_24_inner_macOut = ($signed(_zz__zz__1_24_inner_macOut) + $signed(_zz__zz__1_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_24_inner_activation <= 8'h00;
      _1_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_24_inner_activation <= io_addInput;
      end else begin
        _1_24_inner_macOut <= _zz__1_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_55 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_23_inner_macOut;
  wire       [15:0]   _zz__zz__1_23_inner_macOut_1;
  wire       [15:0]   _zz__1_23_inner_macOut_1;
  wire       [15:0]   _zz__1_23_inner_macOut_2;
  reg        [7:0]    _1_23_inner_activation;
  reg        [7:0]    _1_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_23_inner_macOut;

  assign _zz__zz__1_23_inner_macOut = ($signed(io_mulInput) * $signed(_1_23_inner_activation));
  assign _zz__zz__1_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_23_inner_macOut)) ? 16'h007f : _zz__1_23_inner_macOut_2);
  assign _zz__1_23_inner_macOut_2 = (($signed(_zz__1_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_23_inner_activation;
    end else begin
      io_macOut = _1_23_inner_macOut;
    end
  end

  assign _zz__1_23_inner_macOut = ($signed(_zz__zz__1_23_inner_macOut) + $signed(_zz__zz__1_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_23_inner_activation <= 8'h00;
      _1_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_23_inner_activation <= io_addInput;
      end else begin
        _1_23_inner_macOut <= _zz__1_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_54 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_22_inner_macOut;
  wire       [15:0]   _zz__zz__1_22_inner_macOut_1;
  wire       [15:0]   _zz__1_22_inner_macOut_1;
  wire       [15:0]   _zz__1_22_inner_macOut_2;
  reg        [7:0]    _1_22_inner_activation;
  reg        [7:0]    _1_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_22_inner_macOut;

  assign _zz__zz__1_22_inner_macOut = ($signed(io_mulInput) * $signed(_1_22_inner_activation));
  assign _zz__zz__1_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_22_inner_macOut)) ? 16'h007f : _zz__1_22_inner_macOut_2);
  assign _zz__1_22_inner_macOut_2 = (($signed(_zz__1_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_22_inner_activation;
    end else begin
      io_macOut = _1_22_inner_macOut;
    end
  end

  assign _zz__1_22_inner_macOut = ($signed(_zz__zz__1_22_inner_macOut) + $signed(_zz__zz__1_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_22_inner_activation <= 8'h00;
      _1_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_22_inner_activation <= io_addInput;
      end else begin
        _1_22_inner_macOut <= _zz__1_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_53 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_21_inner_macOut;
  wire       [15:0]   _zz__zz__1_21_inner_macOut_1;
  wire       [15:0]   _zz__1_21_inner_macOut_1;
  wire       [15:0]   _zz__1_21_inner_macOut_2;
  reg        [7:0]    _1_21_inner_activation;
  reg        [7:0]    _1_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_21_inner_macOut;

  assign _zz__zz__1_21_inner_macOut = ($signed(io_mulInput) * $signed(_1_21_inner_activation));
  assign _zz__zz__1_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_21_inner_macOut)) ? 16'h007f : _zz__1_21_inner_macOut_2);
  assign _zz__1_21_inner_macOut_2 = (($signed(_zz__1_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_21_inner_activation;
    end else begin
      io_macOut = _1_21_inner_macOut;
    end
  end

  assign _zz__1_21_inner_macOut = ($signed(_zz__zz__1_21_inner_macOut) + $signed(_zz__zz__1_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_21_inner_activation <= 8'h00;
      _1_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_21_inner_activation <= io_addInput;
      end else begin
        _1_21_inner_macOut <= _zz__1_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_52 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_20_inner_macOut;
  wire       [15:0]   _zz__zz__1_20_inner_macOut_1;
  wire       [15:0]   _zz__1_20_inner_macOut_1;
  wire       [15:0]   _zz__1_20_inner_macOut_2;
  reg        [7:0]    _1_20_inner_activation;
  reg        [7:0]    _1_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_20_inner_macOut;

  assign _zz__zz__1_20_inner_macOut = ($signed(io_mulInput) * $signed(_1_20_inner_activation));
  assign _zz__zz__1_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_20_inner_macOut)) ? 16'h007f : _zz__1_20_inner_macOut_2);
  assign _zz__1_20_inner_macOut_2 = (($signed(_zz__1_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_20_inner_activation;
    end else begin
      io_macOut = _1_20_inner_macOut;
    end
  end

  assign _zz__1_20_inner_macOut = ($signed(_zz__zz__1_20_inner_macOut) + $signed(_zz__zz__1_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_20_inner_activation <= 8'h00;
      _1_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_20_inner_activation <= io_addInput;
      end else begin
        _1_20_inner_macOut <= _zz__1_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_51 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_19_inner_macOut;
  wire       [15:0]   _zz__zz__1_19_inner_macOut_1;
  wire       [15:0]   _zz__1_19_inner_macOut_1;
  wire       [15:0]   _zz__1_19_inner_macOut_2;
  reg        [7:0]    _1_19_inner_activation;
  reg        [7:0]    _1_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_19_inner_macOut;

  assign _zz__zz__1_19_inner_macOut = ($signed(io_mulInput) * $signed(_1_19_inner_activation));
  assign _zz__zz__1_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_19_inner_macOut)) ? 16'h007f : _zz__1_19_inner_macOut_2);
  assign _zz__1_19_inner_macOut_2 = (($signed(_zz__1_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_19_inner_activation;
    end else begin
      io_macOut = _1_19_inner_macOut;
    end
  end

  assign _zz__1_19_inner_macOut = ($signed(_zz__zz__1_19_inner_macOut) + $signed(_zz__zz__1_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_19_inner_activation <= 8'h00;
      _1_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_19_inner_activation <= io_addInput;
      end else begin
        _1_19_inner_macOut <= _zz__1_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_50 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_18_inner_macOut;
  wire       [15:0]   _zz__zz__1_18_inner_macOut_1;
  wire       [15:0]   _zz__1_18_inner_macOut_1;
  wire       [15:0]   _zz__1_18_inner_macOut_2;
  reg        [7:0]    _1_18_inner_activation;
  reg        [7:0]    _1_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_18_inner_macOut;

  assign _zz__zz__1_18_inner_macOut = ($signed(io_mulInput) * $signed(_1_18_inner_activation));
  assign _zz__zz__1_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_18_inner_macOut)) ? 16'h007f : _zz__1_18_inner_macOut_2);
  assign _zz__1_18_inner_macOut_2 = (($signed(_zz__1_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_18_inner_activation;
    end else begin
      io_macOut = _1_18_inner_macOut;
    end
  end

  assign _zz__1_18_inner_macOut = ($signed(_zz__zz__1_18_inner_macOut) + $signed(_zz__zz__1_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_18_inner_activation <= 8'h00;
      _1_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_18_inner_activation <= io_addInput;
      end else begin
        _1_18_inner_macOut <= _zz__1_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_49 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_17_inner_macOut;
  wire       [15:0]   _zz__zz__1_17_inner_macOut_1;
  wire       [15:0]   _zz__1_17_inner_macOut_1;
  wire       [15:0]   _zz__1_17_inner_macOut_2;
  reg        [7:0]    _1_17_inner_activation;
  reg        [7:0]    _1_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_17_inner_macOut;

  assign _zz__zz__1_17_inner_macOut = ($signed(io_mulInput) * $signed(_1_17_inner_activation));
  assign _zz__zz__1_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_17_inner_macOut)) ? 16'h007f : _zz__1_17_inner_macOut_2);
  assign _zz__1_17_inner_macOut_2 = (($signed(_zz__1_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_17_inner_activation;
    end else begin
      io_macOut = _1_17_inner_macOut;
    end
  end

  assign _zz__1_17_inner_macOut = ($signed(_zz__zz__1_17_inner_macOut) + $signed(_zz__zz__1_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_17_inner_activation <= 8'h00;
      _1_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_17_inner_activation <= io_addInput;
      end else begin
        _1_17_inner_macOut <= _zz__1_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_48 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_16_inner_macOut;
  wire       [15:0]   _zz__zz__1_16_inner_macOut_1;
  wire       [15:0]   _zz__1_16_inner_macOut_1;
  wire       [15:0]   _zz__1_16_inner_macOut_2;
  reg        [7:0]    _1_16_inner_activation;
  reg        [7:0]    _1_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_16_inner_macOut;

  assign _zz__zz__1_16_inner_macOut = ($signed(io_mulInput) * $signed(_1_16_inner_activation));
  assign _zz__zz__1_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_16_inner_macOut)) ? 16'h007f : _zz__1_16_inner_macOut_2);
  assign _zz__1_16_inner_macOut_2 = (($signed(_zz__1_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_16_inner_activation;
    end else begin
      io_macOut = _1_16_inner_macOut;
    end
  end

  assign _zz__1_16_inner_macOut = ($signed(_zz__zz__1_16_inner_macOut) + $signed(_zz__zz__1_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_16_inner_activation <= 8'h00;
      _1_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_16_inner_activation <= io_addInput;
      end else begin
        _1_16_inner_macOut <= _zz__1_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_47 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_15_inner_macOut;
  wire       [15:0]   _zz__zz__1_15_inner_macOut_1;
  wire       [15:0]   _zz__1_15_inner_macOut_1;
  wire       [15:0]   _zz__1_15_inner_macOut_2;
  reg        [7:0]    _1_15_inner_activation;
  reg        [7:0]    _1_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_15_inner_macOut;

  assign _zz__zz__1_15_inner_macOut = ($signed(io_mulInput) * $signed(_1_15_inner_activation));
  assign _zz__zz__1_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_15_inner_macOut)) ? 16'h007f : _zz__1_15_inner_macOut_2);
  assign _zz__1_15_inner_macOut_2 = (($signed(_zz__1_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_15_inner_activation;
    end else begin
      io_macOut = _1_15_inner_macOut;
    end
  end

  assign _zz__1_15_inner_macOut = ($signed(_zz__zz__1_15_inner_macOut) + $signed(_zz__zz__1_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_15_inner_activation <= 8'h00;
      _1_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_15_inner_activation <= io_addInput;
      end else begin
        _1_15_inner_macOut <= _zz__1_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_46 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_14_inner_macOut;
  wire       [15:0]   _zz__zz__1_14_inner_macOut_1;
  wire       [15:0]   _zz__1_14_inner_macOut_1;
  wire       [15:0]   _zz__1_14_inner_macOut_2;
  reg        [7:0]    _1_14_inner_activation;
  reg        [7:0]    _1_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_14_inner_macOut;

  assign _zz__zz__1_14_inner_macOut = ($signed(io_mulInput) * $signed(_1_14_inner_activation));
  assign _zz__zz__1_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_14_inner_macOut)) ? 16'h007f : _zz__1_14_inner_macOut_2);
  assign _zz__1_14_inner_macOut_2 = (($signed(_zz__1_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_14_inner_activation;
    end else begin
      io_macOut = _1_14_inner_macOut;
    end
  end

  assign _zz__1_14_inner_macOut = ($signed(_zz__zz__1_14_inner_macOut) + $signed(_zz__zz__1_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_14_inner_activation <= 8'h00;
      _1_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_14_inner_activation <= io_addInput;
      end else begin
        _1_14_inner_macOut <= _zz__1_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_45 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_13_inner_macOut;
  wire       [15:0]   _zz__zz__1_13_inner_macOut_1;
  wire       [15:0]   _zz__1_13_inner_macOut_1;
  wire       [15:0]   _zz__1_13_inner_macOut_2;
  reg        [7:0]    _1_13_inner_activation;
  reg        [7:0]    _1_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_13_inner_macOut;

  assign _zz__zz__1_13_inner_macOut = ($signed(io_mulInput) * $signed(_1_13_inner_activation));
  assign _zz__zz__1_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_13_inner_macOut)) ? 16'h007f : _zz__1_13_inner_macOut_2);
  assign _zz__1_13_inner_macOut_2 = (($signed(_zz__1_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_13_inner_activation;
    end else begin
      io_macOut = _1_13_inner_macOut;
    end
  end

  assign _zz__1_13_inner_macOut = ($signed(_zz__zz__1_13_inner_macOut) + $signed(_zz__zz__1_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_13_inner_activation <= 8'h00;
      _1_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_13_inner_activation <= io_addInput;
      end else begin
        _1_13_inner_macOut <= _zz__1_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_44 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_12_inner_macOut;
  wire       [15:0]   _zz__zz__1_12_inner_macOut_1;
  wire       [15:0]   _zz__1_12_inner_macOut_1;
  wire       [15:0]   _zz__1_12_inner_macOut_2;
  reg        [7:0]    _1_12_inner_activation;
  reg        [7:0]    _1_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_12_inner_macOut;

  assign _zz__zz__1_12_inner_macOut = ($signed(io_mulInput) * $signed(_1_12_inner_activation));
  assign _zz__zz__1_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_12_inner_macOut)) ? 16'h007f : _zz__1_12_inner_macOut_2);
  assign _zz__1_12_inner_macOut_2 = (($signed(_zz__1_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_12_inner_activation;
    end else begin
      io_macOut = _1_12_inner_macOut;
    end
  end

  assign _zz__1_12_inner_macOut = ($signed(_zz__zz__1_12_inner_macOut) + $signed(_zz__zz__1_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_12_inner_activation <= 8'h00;
      _1_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_12_inner_activation <= io_addInput;
      end else begin
        _1_12_inner_macOut <= _zz__1_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_43 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_11_inner_macOut;
  wire       [15:0]   _zz__zz__1_11_inner_macOut_1;
  wire       [15:0]   _zz__1_11_inner_macOut_1;
  wire       [15:0]   _zz__1_11_inner_macOut_2;
  reg        [7:0]    _1_11_inner_activation;
  reg        [7:0]    _1_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_11_inner_macOut;

  assign _zz__zz__1_11_inner_macOut = ($signed(io_mulInput) * $signed(_1_11_inner_activation));
  assign _zz__zz__1_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_11_inner_macOut)) ? 16'h007f : _zz__1_11_inner_macOut_2);
  assign _zz__1_11_inner_macOut_2 = (($signed(_zz__1_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_11_inner_activation;
    end else begin
      io_macOut = _1_11_inner_macOut;
    end
  end

  assign _zz__1_11_inner_macOut = ($signed(_zz__zz__1_11_inner_macOut) + $signed(_zz__zz__1_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_11_inner_activation <= 8'h00;
      _1_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_11_inner_activation <= io_addInput;
      end else begin
        _1_11_inner_macOut <= _zz__1_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_42 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_10_inner_macOut;
  wire       [15:0]   _zz__zz__1_10_inner_macOut_1;
  wire       [15:0]   _zz__1_10_inner_macOut_1;
  wire       [15:0]   _zz__1_10_inner_macOut_2;
  reg        [7:0]    _1_10_inner_activation;
  reg        [7:0]    _1_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_10_inner_macOut;

  assign _zz__zz__1_10_inner_macOut = ($signed(io_mulInput) * $signed(_1_10_inner_activation));
  assign _zz__zz__1_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_10_inner_macOut)) ? 16'h007f : _zz__1_10_inner_macOut_2);
  assign _zz__1_10_inner_macOut_2 = (($signed(_zz__1_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_10_inner_activation;
    end else begin
      io_macOut = _1_10_inner_macOut;
    end
  end

  assign _zz__1_10_inner_macOut = ($signed(_zz__zz__1_10_inner_macOut) + $signed(_zz__zz__1_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_10_inner_activation <= 8'h00;
      _1_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_10_inner_activation <= io_addInput;
      end else begin
        _1_10_inner_macOut <= _zz__1_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_41 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_9_inner_macOut;
  wire       [15:0]   _zz__zz__1_9_inner_macOut_1;
  wire       [15:0]   _zz__1_9_inner_macOut_1;
  wire       [15:0]   _zz__1_9_inner_macOut_2;
  reg        [7:0]    _1_9_inner_activation;
  reg        [7:0]    _1_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_9_inner_macOut;

  assign _zz__zz__1_9_inner_macOut = ($signed(io_mulInput) * $signed(_1_9_inner_activation));
  assign _zz__zz__1_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_9_inner_macOut)) ? 16'h007f : _zz__1_9_inner_macOut_2);
  assign _zz__1_9_inner_macOut_2 = (($signed(_zz__1_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_9_inner_activation;
    end else begin
      io_macOut = _1_9_inner_macOut;
    end
  end

  assign _zz__1_9_inner_macOut = ($signed(_zz__zz__1_9_inner_macOut) + $signed(_zz__zz__1_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_9_inner_activation <= 8'h00;
      _1_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_9_inner_activation <= io_addInput;
      end else begin
        _1_9_inner_macOut <= _zz__1_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_40 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_8_inner_macOut;
  wire       [15:0]   _zz__zz__1_8_inner_macOut_1;
  wire       [15:0]   _zz__1_8_inner_macOut_1;
  wire       [15:0]   _zz__1_8_inner_macOut_2;
  reg        [7:0]    _1_8_inner_activation;
  reg        [7:0]    _1_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_8_inner_macOut;

  assign _zz__zz__1_8_inner_macOut = ($signed(io_mulInput) * $signed(_1_8_inner_activation));
  assign _zz__zz__1_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_8_inner_macOut)) ? 16'h007f : _zz__1_8_inner_macOut_2);
  assign _zz__1_8_inner_macOut_2 = (($signed(_zz__1_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_8_inner_activation;
    end else begin
      io_macOut = _1_8_inner_macOut;
    end
  end

  assign _zz__1_8_inner_macOut = ($signed(_zz__zz__1_8_inner_macOut) + $signed(_zz__zz__1_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_8_inner_activation <= 8'h00;
      _1_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_8_inner_activation <= io_addInput;
      end else begin
        _1_8_inner_macOut <= _zz__1_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_39 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_7_inner_macOut;
  wire       [15:0]   _zz__zz__1_7_inner_macOut_1;
  wire       [15:0]   _zz__1_7_inner_macOut_1;
  wire       [15:0]   _zz__1_7_inner_macOut_2;
  reg        [7:0]    _1_7_inner_activation;
  reg        [7:0]    _1_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_7_inner_macOut;

  assign _zz__zz__1_7_inner_macOut = ($signed(io_mulInput) * $signed(_1_7_inner_activation));
  assign _zz__zz__1_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_7_inner_macOut)) ? 16'h007f : _zz__1_7_inner_macOut_2);
  assign _zz__1_7_inner_macOut_2 = (($signed(_zz__1_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_7_inner_activation;
    end else begin
      io_macOut = _1_7_inner_macOut;
    end
  end

  assign _zz__1_7_inner_macOut = ($signed(_zz__zz__1_7_inner_macOut) + $signed(_zz__zz__1_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_7_inner_activation <= 8'h00;
      _1_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_7_inner_activation <= io_addInput;
      end else begin
        _1_7_inner_macOut <= _zz__1_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_38 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_6_inner_macOut;
  wire       [15:0]   _zz__zz__1_6_inner_macOut_1;
  wire       [15:0]   _zz__1_6_inner_macOut_1;
  wire       [15:0]   _zz__1_6_inner_macOut_2;
  reg        [7:0]    _1_6_inner_activation;
  reg        [7:0]    _1_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_6_inner_macOut;

  assign _zz__zz__1_6_inner_macOut = ($signed(io_mulInput) * $signed(_1_6_inner_activation));
  assign _zz__zz__1_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_6_inner_macOut)) ? 16'h007f : _zz__1_6_inner_macOut_2);
  assign _zz__1_6_inner_macOut_2 = (($signed(_zz__1_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_6_inner_activation;
    end else begin
      io_macOut = _1_6_inner_macOut;
    end
  end

  assign _zz__1_6_inner_macOut = ($signed(_zz__zz__1_6_inner_macOut) + $signed(_zz__zz__1_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_6_inner_activation <= 8'h00;
      _1_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_6_inner_activation <= io_addInput;
      end else begin
        _1_6_inner_macOut <= _zz__1_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_37 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_5_inner_macOut;
  wire       [15:0]   _zz__zz__1_5_inner_macOut_1;
  wire       [15:0]   _zz__1_5_inner_macOut_1;
  wire       [15:0]   _zz__1_5_inner_macOut_2;
  reg        [7:0]    _1_5_inner_activation;
  reg        [7:0]    _1_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_5_inner_macOut;

  assign _zz__zz__1_5_inner_macOut = ($signed(io_mulInput) * $signed(_1_5_inner_activation));
  assign _zz__zz__1_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_5_inner_macOut)) ? 16'h007f : _zz__1_5_inner_macOut_2);
  assign _zz__1_5_inner_macOut_2 = (($signed(_zz__1_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_5_inner_activation;
    end else begin
      io_macOut = _1_5_inner_macOut;
    end
  end

  assign _zz__1_5_inner_macOut = ($signed(_zz__zz__1_5_inner_macOut) + $signed(_zz__zz__1_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_5_inner_activation <= 8'h00;
      _1_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_5_inner_activation <= io_addInput;
      end else begin
        _1_5_inner_macOut <= _zz__1_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_36 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_4_inner_macOut;
  wire       [15:0]   _zz__zz__1_4_inner_macOut_1;
  wire       [15:0]   _zz__1_4_inner_macOut_1;
  wire       [15:0]   _zz__1_4_inner_macOut_2;
  reg        [7:0]    _1_4_inner_activation;
  reg        [7:0]    _1_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_4_inner_macOut;

  assign _zz__zz__1_4_inner_macOut = ($signed(io_mulInput) * $signed(_1_4_inner_activation));
  assign _zz__zz__1_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_4_inner_macOut)) ? 16'h007f : _zz__1_4_inner_macOut_2);
  assign _zz__1_4_inner_macOut_2 = (($signed(_zz__1_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_4_inner_activation;
    end else begin
      io_macOut = _1_4_inner_macOut;
    end
  end

  assign _zz__1_4_inner_macOut = ($signed(_zz__zz__1_4_inner_macOut) + $signed(_zz__zz__1_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_4_inner_activation <= 8'h00;
      _1_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_4_inner_activation <= io_addInput;
      end else begin
        _1_4_inner_macOut <= _zz__1_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_35 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_3_inner_macOut;
  wire       [15:0]   _zz__zz__1_3_inner_macOut_1;
  wire       [15:0]   _zz__1_3_inner_macOut_1;
  wire       [15:0]   _zz__1_3_inner_macOut_2;
  reg        [7:0]    _1_3_inner_activation;
  reg        [7:0]    _1_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_3_inner_macOut;

  assign _zz__zz__1_3_inner_macOut = ($signed(io_mulInput) * $signed(_1_3_inner_activation));
  assign _zz__zz__1_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_3_inner_macOut)) ? 16'h007f : _zz__1_3_inner_macOut_2);
  assign _zz__1_3_inner_macOut_2 = (($signed(_zz__1_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_3_inner_activation;
    end else begin
      io_macOut = _1_3_inner_macOut;
    end
  end

  assign _zz__1_3_inner_macOut = ($signed(_zz__zz__1_3_inner_macOut) + $signed(_zz__zz__1_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_3_inner_activation <= 8'h00;
      _1_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_3_inner_activation <= io_addInput;
      end else begin
        _1_3_inner_macOut <= _zz__1_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_34 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_2_inner_macOut;
  wire       [15:0]   _zz__zz__1_2_inner_macOut_1;
  wire       [15:0]   _zz__1_2_inner_macOut_1;
  wire       [15:0]   _zz__1_2_inner_macOut_2;
  reg        [7:0]    _1_2_inner_activation;
  reg        [7:0]    _1_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_2_inner_macOut;

  assign _zz__zz__1_2_inner_macOut = ($signed(io_mulInput) * $signed(_1_2_inner_activation));
  assign _zz__zz__1_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_2_inner_macOut)) ? 16'h007f : _zz__1_2_inner_macOut_2);
  assign _zz__1_2_inner_macOut_2 = (($signed(_zz__1_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_2_inner_activation;
    end else begin
      io_macOut = _1_2_inner_macOut;
    end
  end

  assign _zz__1_2_inner_macOut = ($signed(_zz__zz__1_2_inner_macOut) + $signed(_zz__zz__1_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_2_inner_activation <= 8'h00;
      _1_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_2_inner_activation <= io_addInput;
      end else begin
        _1_2_inner_macOut <= _zz__1_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_33 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_1_inner_macOut;
  wire       [15:0]   _zz__zz__1_1_inner_macOut_1;
  wire       [15:0]   _zz__1_1_inner_macOut_1;
  wire       [15:0]   _zz__1_1_inner_macOut_2;
  reg        [7:0]    _1_1_inner_activation;
  reg        [7:0]    _1_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_1_inner_macOut;

  assign _zz__zz__1_1_inner_macOut = ($signed(io_mulInput) * $signed(_1_1_inner_activation));
  assign _zz__zz__1_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_1_inner_macOut)) ? 16'h007f : _zz__1_1_inner_macOut_2);
  assign _zz__1_1_inner_macOut_2 = (($signed(_zz__1_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_1_inner_activation;
    end else begin
      io_macOut = _1_1_inner_macOut;
    end
  end

  assign _zz__1_1_inner_macOut = ($signed(_zz__zz__1_1_inner_macOut) + $signed(_zz__zz__1_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_1_inner_activation <= 8'h00;
      _1_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_1_inner_activation <= io_addInput;
      end else begin
        _1_1_inner_macOut <= _zz__1_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_32 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__1_0_inner_macOut;
  wire       [15:0]   _zz__zz__1_0_inner_macOut_1;
  wire       [15:0]   _zz__1_0_inner_macOut_1;
  wire       [15:0]   _zz__1_0_inner_macOut_2;
  reg        [7:0]    _1_0_inner_activation;
  reg        [7:0]    _1_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__1_0_inner_macOut;

  assign _zz__zz__1_0_inner_macOut = ($signed(io_mulInput) * $signed(_1_0_inner_activation));
  assign _zz__zz__1_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__1_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__1_0_inner_macOut)) ? 16'h007f : _zz__1_0_inner_macOut_2);
  assign _zz__1_0_inner_macOut_2 = (($signed(_zz__1_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__1_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _1_0_inner_activation;
    end else begin
      io_macOut = _1_0_inner_macOut;
    end
  end

  assign _zz__1_0_inner_macOut = ($signed(_zz__zz__1_0_inner_macOut) + $signed(_zz__zz__1_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _1_0_inner_activation <= 8'h00;
      _1_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _1_0_inner_activation <= io_addInput;
      end else begin
        _1_0_inner_macOut <= _zz__1_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_31 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_31_inner_macOut;
  wire       [15:0]   _zz__zz__0_31_inner_macOut_1;
  wire       [15:0]   _zz__0_31_inner_macOut_1;
  wire       [15:0]   _zz__0_31_inner_macOut_2;
  reg        [7:0]    _0_31_inner_activation;
  reg        [7:0]    _0_31_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_31_inner_macOut;

  assign _zz__zz__0_31_inner_macOut = ($signed(io_mulInput) * $signed(_0_31_inner_activation));
  assign _zz__zz__0_31_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_31_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_31_inner_macOut)) ? 16'h007f : _zz__0_31_inner_macOut_2);
  assign _zz__0_31_inner_macOut_2 = (($signed(_zz__0_31_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_31_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_31_inner_activation;
    end else begin
      io_macOut = _0_31_inner_macOut;
    end
  end

  assign _zz__0_31_inner_macOut = ($signed(_zz__zz__0_31_inner_macOut) + $signed(_zz__zz__0_31_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_31_inner_activation <= 8'h00;
      _0_31_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_31_inner_activation <= io_addInput;
      end else begin
        _0_31_inner_macOut <= _zz__0_31_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_30 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_30_inner_macOut;
  wire       [15:0]   _zz__zz__0_30_inner_macOut_1;
  wire       [15:0]   _zz__0_30_inner_macOut_1;
  wire       [15:0]   _zz__0_30_inner_macOut_2;
  reg        [7:0]    _0_30_inner_activation;
  reg        [7:0]    _0_30_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_30_inner_macOut;

  assign _zz__zz__0_30_inner_macOut = ($signed(io_mulInput) * $signed(_0_30_inner_activation));
  assign _zz__zz__0_30_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_30_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_30_inner_macOut)) ? 16'h007f : _zz__0_30_inner_macOut_2);
  assign _zz__0_30_inner_macOut_2 = (($signed(_zz__0_30_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_30_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_30_inner_activation;
    end else begin
      io_macOut = _0_30_inner_macOut;
    end
  end

  assign _zz__0_30_inner_macOut = ($signed(_zz__zz__0_30_inner_macOut) + $signed(_zz__zz__0_30_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_30_inner_activation <= 8'h00;
      _0_30_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_30_inner_activation <= io_addInput;
      end else begin
        _0_30_inner_macOut <= _zz__0_30_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_29 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_29_inner_macOut;
  wire       [15:0]   _zz__zz__0_29_inner_macOut_1;
  wire       [15:0]   _zz__0_29_inner_macOut_1;
  wire       [15:0]   _zz__0_29_inner_macOut_2;
  reg        [7:0]    _0_29_inner_activation;
  reg        [7:0]    _0_29_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_29_inner_macOut;

  assign _zz__zz__0_29_inner_macOut = ($signed(io_mulInput) * $signed(_0_29_inner_activation));
  assign _zz__zz__0_29_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_29_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_29_inner_macOut)) ? 16'h007f : _zz__0_29_inner_macOut_2);
  assign _zz__0_29_inner_macOut_2 = (($signed(_zz__0_29_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_29_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_29_inner_activation;
    end else begin
      io_macOut = _0_29_inner_macOut;
    end
  end

  assign _zz__0_29_inner_macOut = ($signed(_zz__zz__0_29_inner_macOut) + $signed(_zz__zz__0_29_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_29_inner_activation <= 8'h00;
      _0_29_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_29_inner_activation <= io_addInput;
      end else begin
        _0_29_inner_macOut <= _zz__0_29_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_28 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_28_inner_macOut;
  wire       [15:0]   _zz__zz__0_28_inner_macOut_1;
  wire       [15:0]   _zz__0_28_inner_macOut_1;
  wire       [15:0]   _zz__0_28_inner_macOut_2;
  reg        [7:0]    _0_28_inner_activation;
  reg        [7:0]    _0_28_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_28_inner_macOut;

  assign _zz__zz__0_28_inner_macOut = ($signed(io_mulInput) * $signed(_0_28_inner_activation));
  assign _zz__zz__0_28_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_28_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_28_inner_macOut)) ? 16'h007f : _zz__0_28_inner_macOut_2);
  assign _zz__0_28_inner_macOut_2 = (($signed(_zz__0_28_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_28_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_28_inner_activation;
    end else begin
      io_macOut = _0_28_inner_macOut;
    end
  end

  assign _zz__0_28_inner_macOut = ($signed(_zz__zz__0_28_inner_macOut) + $signed(_zz__zz__0_28_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_28_inner_activation <= 8'h00;
      _0_28_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_28_inner_activation <= io_addInput;
      end else begin
        _0_28_inner_macOut <= _zz__0_28_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_27 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_27_inner_macOut;
  wire       [15:0]   _zz__zz__0_27_inner_macOut_1;
  wire       [15:0]   _zz__0_27_inner_macOut_1;
  wire       [15:0]   _zz__0_27_inner_macOut_2;
  reg        [7:0]    _0_27_inner_activation;
  reg        [7:0]    _0_27_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_27_inner_macOut;

  assign _zz__zz__0_27_inner_macOut = ($signed(io_mulInput) * $signed(_0_27_inner_activation));
  assign _zz__zz__0_27_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_27_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_27_inner_macOut)) ? 16'h007f : _zz__0_27_inner_macOut_2);
  assign _zz__0_27_inner_macOut_2 = (($signed(_zz__0_27_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_27_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_27_inner_activation;
    end else begin
      io_macOut = _0_27_inner_macOut;
    end
  end

  assign _zz__0_27_inner_macOut = ($signed(_zz__zz__0_27_inner_macOut) + $signed(_zz__zz__0_27_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_27_inner_activation <= 8'h00;
      _0_27_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_27_inner_activation <= io_addInput;
      end else begin
        _0_27_inner_macOut <= _zz__0_27_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_26 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_26_inner_macOut;
  wire       [15:0]   _zz__zz__0_26_inner_macOut_1;
  wire       [15:0]   _zz__0_26_inner_macOut_1;
  wire       [15:0]   _zz__0_26_inner_macOut_2;
  reg        [7:0]    _0_26_inner_activation;
  reg        [7:0]    _0_26_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_26_inner_macOut;

  assign _zz__zz__0_26_inner_macOut = ($signed(io_mulInput) * $signed(_0_26_inner_activation));
  assign _zz__zz__0_26_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_26_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_26_inner_macOut)) ? 16'h007f : _zz__0_26_inner_macOut_2);
  assign _zz__0_26_inner_macOut_2 = (($signed(_zz__0_26_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_26_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_26_inner_activation;
    end else begin
      io_macOut = _0_26_inner_macOut;
    end
  end

  assign _zz__0_26_inner_macOut = ($signed(_zz__zz__0_26_inner_macOut) + $signed(_zz__zz__0_26_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_26_inner_activation <= 8'h00;
      _0_26_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_26_inner_activation <= io_addInput;
      end else begin
        _0_26_inner_macOut <= _zz__0_26_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_25 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_25_inner_macOut;
  wire       [15:0]   _zz__zz__0_25_inner_macOut_1;
  wire       [15:0]   _zz__0_25_inner_macOut_1;
  wire       [15:0]   _zz__0_25_inner_macOut_2;
  reg        [7:0]    _0_25_inner_activation;
  reg        [7:0]    _0_25_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_25_inner_macOut;

  assign _zz__zz__0_25_inner_macOut = ($signed(io_mulInput) * $signed(_0_25_inner_activation));
  assign _zz__zz__0_25_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_25_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_25_inner_macOut)) ? 16'h007f : _zz__0_25_inner_macOut_2);
  assign _zz__0_25_inner_macOut_2 = (($signed(_zz__0_25_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_25_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_25_inner_activation;
    end else begin
      io_macOut = _0_25_inner_macOut;
    end
  end

  assign _zz__0_25_inner_macOut = ($signed(_zz__zz__0_25_inner_macOut) + $signed(_zz__zz__0_25_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_25_inner_activation <= 8'h00;
      _0_25_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_25_inner_activation <= io_addInput;
      end else begin
        _0_25_inner_macOut <= _zz__0_25_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_24 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_24_inner_macOut;
  wire       [15:0]   _zz__zz__0_24_inner_macOut_1;
  wire       [15:0]   _zz__0_24_inner_macOut_1;
  wire       [15:0]   _zz__0_24_inner_macOut_2;
  reg        [7:0]    _0_24_inner_activation;
  reg        [7:0]    _0_24_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_24_inner_macOut;

  assign _zz__zz__0_24_inner_macOut = ($signed(io_mulInput) * $signed(_0_24_inner_activation));
  assign _zz__zz__0_24_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_24_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_24_inner_macOut)) ? 16'h007f : _zz__0_24_inner_macOut_2);
  assign _zz__0_24_inner_macOut_2 = (($signed(_zz__0_24_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_24_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_24_inner_activation;
    end else begin
      io_macOut = _0_24_inner_macOut;
    end
  end

  assign _zz__0_24_inner_macOut = ($signed(_zz__zz__0_24_inner_macOut) + $signed(_zz__zz__0_24_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_24_inner_activation <= 8'h00;
      _0_24_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_24_inner_activation <= io_addInput;
      end else begin
        _0_24_inner_macOut <= _zz__0_24_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_23 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_23_inner_macOut;
  wire       [15:0]   _zz__zz__0_23_inner_macOut_1;
  wire       [15:0]   _zz__0_23_inner_macOut_1;
  wire       [15:0]   _zz__0_23_inner_macOut_2;
  reg        [7:0]    _0_23_inner_activation;
  reg        [7:0]    _0_23_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_23_inner_macOut;

  assign _zz__zz__0_23_inner_macOut = ($signed(io_mulInput) * $signed(_0_23_inner_activation));
  assign _zz__zz__0_23_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_23_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_23_inner_macOut)) ? 16'h007f : _zz__0_23_inner_macOut_2);
  assign _zz__0_23_inner_macOut_2 = (($signed(_zz__0_23_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_23_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_23_inner_activation;
    end else begin
      io_macOut = _0_23_inner_macOut;
    end
  end

  assign _zz__0_23_inner_macOut = ($signed(_zz__zz__0_23_inner_macOut) + $signed(_zz__zz__0_23_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_23_inner_activation <= 8'h00;
      _0_23_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_23_inner_activation <= io_addInput;
      end else begin
        _0_23_inner_macOut <= _zz__0_23_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_22 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_22_inner_macOut;
  wire       [15:0]   _zz__zz__0_22_inner_macOut_1;
  wire       [15:0]   _zz__0_22_inner_macOut_1;
  wire       [15:0]   _zz__0_22_inner_macOut_2;
  reg        [7:0]    _0_22_inner_activation;
  reg        [7:0]    _0_22_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_22_inner_macOut;

  assign _zz__zz__0_22_inner_macOut = ($signed(io_mulInput) * $signed(_0_22_inner_activation));
  assign _zz__zz__0_22_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_22_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_22_inner_macOut)) ? 16'h007f : _zz__0_22_inner_macOut_2);
  assign _zz__0_22_inner_macOut_2 = (($signed(_zz__0_22_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_22_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_22_inner_activation;
    end else begin
      io_macOut = _0_22_inner_macOut;
    end
  end

  assign _zz__0_22_inner_macOut = ($signed(_zz__zz__0_22_inner_macOut) + $signed(_zz__zz__0_22_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_22_inner_activation <= 8'h00;
      _0_22_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_22_inner_activation <= io_addInput;
      end else begin
        _0_22_inner_macOut <= _zz__0_22_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_21 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_21_inner_macOut;
  wire       [15:0]   _zz__zz__0_21_inner_macOut_1;
  wire       [15:0]   _zz__0_21_inner_macOut_1;
  wire       [15:0]   _zz__0_21_inner_macOut_2;
  reg        [7:0]    _0_21_inner_activation;
  reg        [7:0]    _0_21_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_21_inner_macOut;

  assign _zz__zz__0_21_inner_macOut = ($signed(io_mulInput) * $signed(_0_21_inner_activation));
  assign _zz__zz__0_21_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_21_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_21_inner_macOut)) ? 16'h007f : _zz__0_21_inner_macOut_2);
  assign _zz__0_21_inner_macOut_2 = (($signed(_zz__0_21_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_21_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_21_inner_activation;
    end else begin
      io_macOut = _0_21_inner_macOut;
    end
  end

  assign _zz__0_21_inner_macOut = ($signed(_zz__zz__0_21_inner_macOut) + $signed(_zz__zz__0_21_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_21_inner_activation <= 8'h00;
      _0_21_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_21_inner_activation <= io_addInput;
      end else begin
        _0_21_inner_macOut <= _zz__0_21_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_20 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_20_inner_macOut;
  wire       [15:0]   _zz__zz__0_20_inner_macOut_1;
  wire       [15:0]   _zz__0_20_inner_macOut_1;
  wire       [15:0]   _zz__0_20_inner_macOut_2;
  reg        [7:0]    _0_20_inner_activation;
  reg        [7:0]    _0_20_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_20_inner_macOut;

  assign _zz__zz__0_20_inner_macOut = ($signed(io_mulInput) * $signed(_0_20_inner_activation));
  assign _zz__zz__0_20_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_20_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_20_inner_macOut)) ? 16'h007f : _zz__0_20_inner_macOut_2);
  assign _zz__0_20_inner_macOut_2 = (($signed(_zz__0_20_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_20_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_20_inner_activation;
    end else begin
      io_macOut = _0_20_inner_macOut;
    end
  end

  assign _zz__0_20_inner_macOut = ($signed(_zz__zz__0_20_inner_macOut) + $signed(_zz__zz__0_20_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_20_inner_activation <= 8'h00;
      _0_20_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_20_inner_activation <= io_addInput;
      end else begin
        _0_20_inner_macOut <= _zz__0_20_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_19 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_19_inner_macOut;
  wire       [15:0]   _zz__zz__0_19_inner_macOut_1;
  wire       [15:0]   _zz__0_19_inner_macOut_1;
  wire       [15:0]   _zz__0_19_inner_macOut_2;
  reg        [7:0]    _0_19_inner_activation;
  reg        [7:0]    _0_19_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_19_inner_macOut;

  assign _zz__zz__0_19_inner_macOut = ($signed(io_mulInput) * $signed(_0_19_inner_activation));
  assign _zz__zz__0_19_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_19_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_19_inner_macOut)) ? 16'h007f : _zz__0_19_inner_macOut_2);
  assign _zz__0_19_inner_macOut_2 = (($signed(_zz__0_19_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_19_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_19_inner_activation;
    end else begin
      io_macOut = _0_19_inner_macOut;
    end
  end

  assign _zz__0_19_inner_macOut = ($signed(_zz__zz__0_19_inner_macOut) + $signed(_zz__zz__0_19_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_19_inner_activation <= 8'h00;
      _0_19_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_19_inner_activation <= io_addInput;
      end else begin
        _0_19_inner_macOut <= _zz__0_19_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_18 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_18_inner_macOut;
  wire       [15:0]   _zz__zz__0_18_inner_macOut_1;
  wire       [15:0]   _zz__0_18_inner_macOut_1;
  wire       [15:0]   _zz__0_18_inner_macOut_2;
  reg        [7:0]    _0_18_inner_activation;
  reg        [7:0]    _0_18_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_18_inner_macOut;

  assign _zz__zz__0_18_inner_macOut = ($signed(io_mulInput) * $signed(_0_18_inner_activation));
  assign _zz__zz__0_18_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_18_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_18_inner_macOut)) ? 16'h007f : _zz__0_18_inner_macOut_2);
  assign _zz__0_18_inner_macOut_2 = (($signed(_zz__0_18_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_18_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_18_inner_activation;
    end else begin
      io_macOut = _0_18_inner_macOut;
    end
  end

  assign _zz__0_18_inner_macOut = ($signed(_zz__zz__0_18_inner_macOut) + $signed(_zz__zz__0_18_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_18_inner_activation <= 8'h00;
      _0_18_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_18_inner_activation <= io_addInput;
      end else begin
        _0_18_inner_macOut <= _zz__0_18_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_17 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_17_inner_macOut;
  wire       [15:0]   _zz__zz__0_17_inner_macOut_1;
  wire       [15:0]   _zz__0_17_inner_macOut_1;
  wire       [15:0]   _zz__0_17_inner_macOut_2;
  reg        [7:0]    _0_17_inner_activation;
  reg        [7:0]    _0_17_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_17_inner_macOut;

  assign _zz__zz__0_17_inner_macOut = ($signed(io_mulInput) * $signed(_0_17_inner_activation));
  assign _zz__zz__0_17_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_17_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_17_inner_macOut)) ? 16'h007f : _zz__0_17_inner_macOut_2);
  assign _zz__0_17_inner_macOut_2 = (($signed(_zz__0_17_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_17_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_17_inner_activation;
    end else begin
      io_macOut = _0_17_inner_macOut;
    end
  end

  assign _zz__0_17_inner_macOut = ($signed(_zz__zz__0_17_inner_macOut) + $signed(_zz__zz__0_17_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_17_inner_activation <= 8'h00;
      _0_17_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_17_inner_activation <= io_addInput;
      end else begin
        _0_17_inner_macOut <= _zz__0_17_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_16 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_16_inner_macOut;
  wire       [15:0]   _zz__zz__0_16_inner_macOut_1;
  wire       [15:0]   _zz__0_16_inner_macOut_1;
  wire       [15:0]   _zz__0_16_inner_macOut_2;
  reg        [7:0]    _0_16_inner_activation;
  reg        [7:0]    _0_16_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_16_inner_macOut;

  assign _zz__zz__0_16_inner_macOut = ($signed(io_mulInput) * $signed(_0_16_inner_activation));
  assign _zz__zz__0_16_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_16_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_16_inner_macOut)) ? 16'h007f : _zz__0_16_inner_macOut_2);
  assign _zz__0_16_inner_macOut_2 = (($signed(_zz__0_16_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_16_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_16_inner_activation;
    end else begin
      io_macOut = _0_16_inner_macOut;
    end
  end

  assign _zz__0_16_inner_macOut = ($signed(_zz__zz__0_16_inner_macOut) + $signed(_zz__zz__0_16_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_16_inner_activation <= 8'h00;
      _0_16_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_16_inner_activation <= io_addInput;
      end else begin
        _0_16_inner_macOut <= _zz__0_16_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_15 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_15_inner_macOut;
  wire       [15:0]   _zz__zz__0_15_inner_macOut_1;
  wire       [15:0]   _zz__0_15_inner_macOut_1;
  wire       [15:0]   _zz__0_15_inner_macOut_2;
  reg        [7:0]    _0_15_inner_activation;
  reg        [7:0]    _0_15_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_15_inner_macOut;

  assign _zz__zz__0_15_inner_macOut = ($signed(io_mulInput) * $signed(_0_15_inner_activation));
  assign _zz__zz__0_15_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_15_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_15_inner_macOut)) ? 16'h007f : _zz__0_15_inner_macOut_2);
  assign _zz__0_15_inner_macOut_2 = (($signed(_zz__0_15_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_15_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_15_inner_activation;
    end else begin
      io_macOut = _0_15_inner_macOut;
    end
  end

  assign _zz__0_15_inner_macOut = ($signed(_zz__zz__0_15_inner_macOut) + $signed(_zz__zz__0_15_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_15_inner_activation <= 8'h00;
      _0_15_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_15_inner_activation <= io_addInput;
      end else begin
        _0_15_inner_macOut <= _zz__0_15_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_14 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_14_inner_macOut;
  wire       [15:0]   _zz__zz__0_14_inner_macOut_1;
  wire       [15:0]   _zz__0_14_inner_macOut_1;
  wire       [15:0]   _zz__0_14_inner_macOut_2;
  reg        [7:0]    _0_14_inner_activation;
  reg        [7:0]    _0_14_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_14_inner_macOut;

  assign _zz__zz__0_14_inner_macOut = ($signed(io_mulInput) * $signed(_0_14_inner_activation));
  assign _zz__zz__0_14_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_14_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_14_inner_macOut)) ? 16'h007f : _zz__0_14_inner_macOut_2);
  assign _zz__0_14_inner_macOut_2 = (($signed(_zz__0_14_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_14_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_14_inner_activation;
    end else begin
      io_macOut = _0_14_inner_macOut;
    end
  end

  assign _zz__0_14_inner_macOut = ($signed(_zz__zz__0_14_inner_macOut) + $signed(_zz__zz__0_14_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_14_inner_activation <= 8'h00;
      _0_14_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_14_inner_activation <= io_addInput;
      end else begin
        _0_14_inner_macOut <= _zz__0_14_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_13 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_13_inner_macOut;
  wire       [15:0]   _zz__zz__0_13_inner_macOut_1;
  wire       [15:0]   _zz__0_13_inner_macOut_1;
  wire       [15:0]   _zz__0_13_inner_macOut_2;
  reg        [7:0]    _0_13_inner_activation;
  reg        [7:0]    _0_13_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_13_inner_macOut;

  assign _zz__zz__0_13_inner_macOut = ($signed(io_mulInput) * $signed(_0_13_inner_activation));
  assign _zz__zz__0_13_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_13_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_13_inner_macOut)) ? 16'h007f : _zz__0_13_inner_macOut_2);
  assign _zz__0_13_inner_macOut_2 = (($signed(_zz__0_13_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_13_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_13_inner_activation;
    end else begin
      io_macOut = _0_13_inner_macOut;
    end
  end

  assign _zz__0_13_inner_macOut = ($signed(_zz__zz__0_13_inner_macOut) + $signed(_zz__zz__0_13_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_13_inner_activation <= 8'h00;
      _0_13_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_13_inner_activation <= io_addInput;
      end else begin
        _0_13_inner_macOut <= _zz__0_13_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_12 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_12_inner_macOut;
  wire       [15:0]   _zz__zz__0_12_inner_macOut_1;
  wire       [15:0]   _zz__0_12_inner_macOut_1;
  wire       [15:0]   _zz__0_12_inner_macOut_2;
  reg        [7:0]    _0_12_inner_activation;
  reg        [7:0]    _0_12_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_12_inner_macOut;

  assign _zz__zz__0_12_inner_macOut = ($signed(io_mulInput) * $signed(_0_12_inner_activation));
  assign _zz__zz__0_12_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_12_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_12_inner_macOut)) ? 16'h007f : _zz__0_12_inner_macOut_2);
  assign _zz__0_12_inner_macOut_2 = (($signed(_zz__0_12_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_12_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_12_inner_activation;
    end else begin
      io_macOut = _0_12_inner_macOut;
    end
  end

  assign _zz__0_12_inner_macOut = ($signed(_zz__zz__0_12_inner_macOut) + $signed(_zz__zz__0_12_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_12_inner_activation <= 8'h00;
      _0_12_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_12_inner_activation <= io_addInput;
      end else begin
        _0_12_inner_macOut <= _zz__0_12_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_11 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_11_inner_macOut;
  wire       [15:0]   _zz__zz__0_11_inner_macOut_1;
  wire       [15:0]   _zz__0_11_inner_macOut_1;
  wire       [15:0]   _zz__0_11_inner_macOut_2;
  reg        [7:0]    _0_11_inner_activation;
  reg        [7:0]    _0_11_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_11_inner_macOut;

  assign _zz__zz__0_11_inner_macOut = ($signed(io_mulInput) * $signed(_0_11_inner_activation));
  assign _zz__zz__0_11_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_11_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_11_inner_macOut)) ? 16'h007f : _zz__0_11_inner_macOut_2);
  assign _zz__0_11_inner_macOut_2 = (($signed(_zz__0_11_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_11_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_11_inner_activation;
    end else begin
      io_macOut = _0_11_inner_macOut;
    end
  end

  assign _zz__0_11_inner_macOut = ($signed(_zz__zz__0_11_inner_macOut) + $signed(_zz__zz__0_11_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_11_inner_activation <= 8'h00;
      _0_11_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_11_inner_activation <= io_addInput;
      end else begin
        _0_11_inner_macOut <= _zz__0_11_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_10 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_10_inner_macOut;
  wire       [15:0]   _zz__zz__0_10_inner_macOut_1;
  wire       [15:0]   _zz__0_10_inner_macOut_1;
  wire       [15:0]   _zz__0_10_inner_macOut_2;
  reg        [7:0]    _0_10_inner_activation;
  reg        [7:0]    _0_10_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_10_inner_macOut;

  assign _zz__zz__0_10_inner_macOut = ($signed(io_mulInput) * $signed(_0_10_inner_activation));
  assign _zz__zz__0_10_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_10_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_10_inner_macOut)) ? 16'h007f : _zz__0_10_inner_macOut_2);
  assign _zz__0_10_inner_macOut_2 = (($signed(_zz__0_10_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_10_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_10_inner_activation;
    end else begin
      io_macOut = _0_10_inner_macOut;
    end
  end

  assign _zz__0_10_inner_macOut = ($signed(_zz__zz__0_10_inner_macOut) + $signed(_zz__zz__0_10_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_10_inner_activation <= 8'h00;
      _0_10_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_10_inner_activation <= io_addInput;
      end else begin
        _0_10_inner_macOut <= _zz__0_10_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_9 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_9_inner_macOut;
  wire       [15:0]   _zz__zz__0_9_inner_macOut_1;
  wire       [15:0]   _zz__0_9_inner_macOut_1;
  wire       [15:0]   _zz__0_9_inner_macOut_2;
  reg        [7:0]    _0_9_inner_activation;
  reg        [7:0]    _0_9_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_9_inner_macOut;

  assign _zz__zz__0_9_inner_macOut = ($signed(io_mulInput) * $signed(_0_9_inner_activation));
  assign _zz__zz__0_9_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_9_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_9_inner_macOut)) ? 16'h007f : _zz__0_9_inner_macOut_2);
  assign _zz__0_9_inner_macOut_2 = (($signed(_zz__0_9_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_9_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_9_inner_activation;
    end else begin
      io_macOut = _0_9_inner_macOut;
    end
  end

  assign _zz__0_9_inner_macOut = ($signed(_zz__zz__0_9_inner_macOut) + $signed(_zz__zz__0_9_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_9_inner_activation <= 8'h00;
      _0_9_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_9_inner_activation <= io_addInput;
      end else begin
        _0_9_inner_macOut <= _zz__0_9_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_8 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_8_inner_macOut;
  wire       [15:0]   _zz__zz__0_8_inner_macOut_1;
  wire       [15:0]   _zz__0_8_inner_macOut_1;
  wire       [15:0]   _zz__0_8_inner_macOut_2;
  reg        [7:0]    _0_8_inner_activation;
  reg        [7:0]    _0_8_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_8_inner_macOut;

  assign _zz__zz__0_8_inner_macOut = ($signed(io_mulInput) * $signed(_0_8_inner_activation));
  assign _zz__zz__0_8_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_8_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_8_inner_macOut)) ? 16'h007f : _zz__0_8_inner_macOut_2);
  assign _zz__0_8_inner_macOut_2 = (($signed(_zz__0_8_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_8_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_8_inner_activation;
    end else begin
      io_macOut = _0_8_inner_macOut;
    end
  end

  assign _zz__0_8_inner_macOut = ($signed(_zz__zz__0_8_inner_macOut) + $signed(_zz__zz__0_8_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_8_inner_activation <= 8'h00;
      _0_8_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_8_inner_activation <= io_addInput;
      end else begin
        _0_8_inner_macOut <= _zz__0_8_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_7 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_7_inner_macOut;
  wire       [15:0]   _zz__zz__0_7_inner_macOut_1;
  wire       [15:0]   _zz__0_7_inner_macOut_1;
  wire       [15:0]   _zz__0_7_inner_macOut_2;
  reg        [7:0]    _0_7_inner_activation;
  reg        [7:0]    _0_7_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_7_inner_macOut;

  assign _zz__zz__0_7_inner_macOut = ($signed(io_mulInput) * $signed(_0_7_inner_activation));
  assign _zz__zz__0_7_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_7_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_7_inner_macOut)) ? 16'h007f : _zz__0_7_inner_macOut_2);
  assign _zz__0_7_inner_macOut_2 = (($signed(_zz__0_7_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_7_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_7_inner_activation;
    end else begin
      io_macOut = _0_7_inner_macOut;
    end
  end

  assign _zz__0_7_inner_macOut = ($signed(_zz__zz__0_7_inner_macOut) + $signed(_zz__zz__0_7_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_7_inner_activation <= 8'h00;
      _0_7_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_7_inner_activation <= io_addInput;
      end else begin
        _0_7_inner_macOut <= _zz__0_7_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_6 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_6_inner_macOut;
  wire       [15:0]   _zz__zz__0_6_inner_macOut_1;
  wire       [15:0]   _zz__0_6_inner_macOut_1;
  wire       [15:0]   _zz__0_6_inner_macOut_2;
  reg        [7:0]    _0_6_inner_activation;
  reg        [7:0]    _0_6_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_6_inner_macOut;

  assign _zz__zz__0_6_inner_macOut = ($signed(io_mulInput) * $signed(_0_6_inner_activation));
  assign _zz__zz__0_6_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_6_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_6_inner_macOut)) ? 16'h007f : _zz__0_6_inner_macOut_2);
  assign _zz__0_6_inner_macOut_2 = (($signed(_zz__0_6_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_6_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_6_inner_activation;
    end else begin
      io_macOut = _0_6_inner_macOut;
    end
  end

  assign _zz__0_6_inner_macOut = ($signed(_zz__zz__0_6_inner_macOut) + $signed(_zz__zz__0_6_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_6_inner_activation <= 8'h00;
      _0_6_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_6_inner_activation <= io_addInput;
      end else begin
        _0_6_inner_macOut <= _zz__0_6_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_5 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_5_inner_macOut;
  wire       [15:0]   _zz__zz__0_5_inner_macOut_1;
  wire       [15:0]   _zz__0_5_inner_macOut_1;
  wire       [15:0]   _zz__0_5_inner_macOut_2;
  reg        [7:0]    _0_5_inner_activation;
  reg        [7:0]    _0_5_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_5_inner_macOut;

  assign _zz__zz__0_5_inner_macOut = ($signed(io_mulInput) * $signed(_0_5_inner_activation));
  assign _zz__zz__0_5_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_5_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_5_inner_macOut)) ? 16'h007f : _zz__0_5_inner_macOut_2);
  assign _zz__0_5_inner_macOut_2 = (($signed(_zz__0_5_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_5_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_5_inner_activation;
    end else begin
      io_macOut = _0_5_inner_macOut;
    end
  end

  assign _zz__0_5_inner_macOut = ($signed(_zz__zz__0_5_inner_macOut) + $signed(_zz__zz__0_5_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_5_inner_activation <= 8'h00;
      _0_5_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_5_inner_activation <= io_addInput;
      end else begin
        _0_5_inner_macOut <= _zz__0_5_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_4 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_4_inner_macOut;
  wire       [15:0]   _zz__zz__0_4_inner_macOut_1;
  wire       [15:0]   _zz__0_4_inner_macOut_1;
  wire       [15:0]   _zz__0_4_inner_macOut_2;
  reg        [7:0]    _0_4_inner_activation;
  reg        [7:0]    _0_4_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_4_inner_macOut;

  assign _zz__zz__0_4_inner_macOut = ($signed(io_mulInput) * $signed(_0_4_inner_activation));
  assign _zz__zz__0_4_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_4_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_4_inner_macOut)) ? 16'h007f : _zz__0_4_inner_macOut_2);
  assign _zz__0_4_inner_macOut_2 = (($signed(_zz__0_4_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_4_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_4_inner_activation;
    end else begin
      io_macOut = _0_4_inner_macOut;
    end
  end

  assign _zz__0_4_inner_macOut = ($signed(_zz__zz__0_4_inner_macOut) + $signed(_zz__zz__0_4_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_4_inner_activation <= 8'h00;
      _0_4_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_4_inner_activation <= io_addInput;
      end else begin
        _0_4_inner_macOut <= _zz__0_4_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_3 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_3_inner_macOut;
  wire       [15:0]   _zz__zz__0_3_inner_macOut_1;
  wire       [15:0]   _zz__0_3_inner_macOut_1;
  wire       [15:0]   _zz__0_3_inner_macOut_2;
  reg        [7:0]    _0_3_inner_activation;
  reg        [7:0]    _0_3_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_3_inner_macOut;

  assign _zz__zz__0_3_inner_macOut = ($signed(io_mulInput) * $signed(_0_3_inner_activation));
  assign _zz__zz__0_3_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_3_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_3_inner_macOut)) ? 16'h007f : _zz__0_3_inner_macOut_2);
  assign _zz__0_3_inner_macOut_2 = (($signed(_zz__0_3_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_3_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_3_inner_activation;
    end else begin
      io_macOut = _0_3_inner_macOut;
    end
  end

  assign _zz__0_3_inner_macOut = ($signed(_zz__zz__0_3_inner_macOut) + $signed(_zz__zz__0_3_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_3_inner_activation <= 8'h00;
      _0_3_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_3_inner_activation <= io_addInput;
      end else begin
        _0_3_inner_macOut <= _zz__0_3_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_2 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_2_inner_macOut;
  wire       [15:0]   _zz__zz__0_2_inner_macOut_1;
  wire       [15:0]   _zz__0_2_inner_macOut_1;
  wire       [15:0]   _zz__0_2_inner_macOut_2;
  reg        [7:0]    _0_2_inner_activation;
  reg        [7:0]    _0_2_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_2_inner_macOut;

  assign _zz__zz__0_2_inner_macOut = ($signed(io_mulInput) * $signed(_0_2_inner_activation));
  assign _zz__zz__0_2_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_2_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_2_inner_macOut)) ? 16'h007f : _zz__0_2_inner_macOut_2);
  assign _zz__0_2_inner_macOut_2 = (($signed(_zz__0_2_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_2_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_2_inner_activation;
    end else begin
      io_macOut = _0_2_inner_macOut;
    end
  end

  assign _zz__0_2_inner_macOut = ($signed(_zz__zz__0_2_inner_macOut) + $signed(_zz__zz__0_2_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_2_inner_activation <= 8'h00;
      _0_2_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_2_inner_activation <= io_addInput;
      end else begin
        _0_2_inner_macOut <= _zz__0_2_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC_1 (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_1_inner_macOut;
  wire       [15:0]   _zz__zz__0_1_inner_macOut_1;
  wire       [15:0]   _zz__0_1_inner_macOut_1;
  wire       [15:0]   _zz__0_1_inner_macOut_2;
  reg        [7:0]    _0_1_inner_activation;
  reg        [7:0]    _0_1_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_1_inner_macOut;

  assign _zz__zz__0_1_inner_macOut = ($signed(io_mulInput) * $signed(_0_1_inner_activation));
  assign _zz__zz__0_1_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_1_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_1_inner_macOut)) ? 16'h007f : _zz__0_1_inner_macOut_2);
  assign _zz__0_1_inner_macOut_2 = (($signed(_zz__0_1_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_1_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_1_inner_activation;
    end else begin
      io_macOut = _0_1_inner_macOut;
    end
  end

  assign _zz__0_1_inner_macOut = ($signed(_zz__zz__0_1_inner_macOut) + $signed(_zz__zz__0_1_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_1_inner_activation <= 8'h00;
      _0_1_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_1_inner_activation <= io_addInput;
      end else begin
        _0_1_inner_macOut <= _zz__0_1_inner_macOut_1[7:0];
      end
    end
  end


endmodule

module MAC (
  input  wire          io_load,
  input  wire [7:0]    io_mulInput,
  input  wire [7:0]    io_addInput,
  output wire [7:0]    io_passthrough,
  output reg  [7:0]    io_macOut,
  input  wire          clk,
  input  wire          reset
);

  wire       [15:0]   _zz__zz__0_0_inner_macOut;
  wire       [15:0]   _zz__zz__0_0_inner_macOut_1;
  wire       [15:0]   _zz__0_0_inner_macOut_1;
  wire       [15:0]   _zz__0_0_inner_macOut_2;
  reg        [7:0]    _0_0_inner_activation;
  reg        [7:0]    _0_0_inner_macOut;
  reg        [7:0]    io_mulInput_regNext;
  wire       [15:0]   _zz__0_0_inner_macOut;

  assign _zz__zz__0_0_inner_macOut = ($signed(io_mulInput) * $signed(_0_0_inner_activation));
  assign _zz__zz__0_0_inner_macOut_1 = {{8{io_addInput[7]}}, io_addInput};
  assign _zz__0_0_inner_macOut_1 = (($signed(16'h007f) < $signed(_zz__0_0_inner_macOut)) ? 16'h007f : _zz__0_0_inner_macOut_2);
  assign _zz__0_0_inner_macOut_2 = (($signed(_zz__0_0_inner_macOut) < $signed(16'hff80)) ? 16'hff80 : _zz__0_0_inner_macOut);
  assign io_passthrough = io_mulInput_regNext;
  always @(*) begin
    if(io_load) begin
      io_macOut = _0_0_inner_activation;
    end else begin
      io_macOut = _0_0_inner_macOut;
    end
  end

  assign _zz__0_0_inner_macOut = ($signed(_zz__zz__0_0_inner_macOut) + $signed(_zz__zz__0_0_inner_macOut_1));
  always @(posedge clk or posedge reset) begin
    if(reset) begin
      _0_0_inner_activation <= 8'h00;
      _0_0_inner_macOut <= 8'h00;
      io_mulInput_regNext <= 8'h00;
    end else begin
      io_mulInput_regNext <= io_mulInput;
      if(io_load) begin
        _0_0_inner_activation <= io_addInput;
      end else begin
        _0_0_inner_macOut <= _zz__0_0_inner_macOut_1[7:0];
      end
    end
  end


endmodule
